library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e0edc287",
    12 => x"86c0c84e",
    13 => x"49e0edc2",
    14 => x"48ccdbc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c6e0",
    19 => x"721e87fd",
    20 => x"121e731e",
    21 => x"ca021148",
    22 => x"dfc34b87",
    23 => x"88739b98",
    24 => x"2687f002",
    25 => x"264a264b",
    26 => x"1e731e4f",
    27 => x"8bc11e72",
    28 => x"1287ca04",
    29 => x"c4021148",
    30 => x"f1028887",
    31 => x"264a2687",
    32 => x"1e4f264b",
    33 => x"1e731e74",
    34 => x"8bc11e72",
    35 => x"1287d004",
    36 => x"ca021148",
    37 => x"dfc34c87",
    38 => x"88749c98",
    39 => x"2687eb02",
    40 => x"264b264a",
    41 => x"1e4f264c",
    42 => x"73814873",
    43 => x"87c502a9",
    44 => x"f6055312",
    45 => x"1e4f2687",
    46 => x"66c44a71",
    47 => x"88c14849",
    48 => x"7158a6c8",
    49 => x"87d40299",
    50 => x"d4ff4812",
    51 => x"66c47808",
    52 => x"88c14849",
    53 => x"7158a6c8",
    54 => x"87ec0599",
    55 => x"711e4f26",
    56 => x"4966c44a",
    57 => x"c888c148",
    58 => x"997158a6",
    59 => x"ff87d602",
    60 => x"ffc348d4",
    61 => x"c4526878",
    62 => x"c1484966",
    63 => x"58a6c888",
    64 => x"ea059971",
    65 => x"1e4f2687",
    66 => x"d4ff1e73",
    67 => x"7bffc34b",
    68 => x"ffc34a6b",
    69 => x"c8496b7b",
    70 => x"c3b17232",
    71 => x"4a6b7bff",
    72 => x"b27131c8",
    73 => x"6b7bffc3",
    74 => x"7232c849",
    75 => x"c44871b1",
    76 => x"264d2687",
    77 => x"264b264c",
    78 => x"5b5e0e4f",
    79 => x"710e5d5c",
    80 => x"4cd4ff4a",
    81 => x"ffc34872",
    82 => x"c27c7098",
    83 => x"05bfccdb",
    84 => x"66d087c8",
    85 => x"d430c948",
    86 => x"66d058a6",
    87 => x"7129d849",
    88 => x"98ffc348",
    89 => x"66d07c70",
    90 => x"7129d049",
    91 => x"98ffc348",
    92 => x"66d07c70",
    93 => x"7129c849",
    94 => x"98ffc348",
    95 => x"66d07c70",
    96 => x"98ffc348",
    97 => x"49727c70",
    98 => x"487129d0",
    99 => x"7098ffc3",
   100 => x"c94b6c7c",
   101 => x"c34dfff0",
   102 => x"d005abff",
   103 => x"7cffc387",
   104 => x"8dc14b6c",
   105 => x"c387c602",
   106 => x"f002abff",
   107 => x"fd487387",
   108 => x"c01e87ff",
   109 => x"48d4ff49",
   110 => x"c178ffc3",
   111 => x"b7c8c381",
   112 => x"87f104a9",
   113 => x"731e4f26",
   114 => x"c487e71e",
   115 => x"c04bdff8",
   116 => x"f0ffc01e",
   117 => x"fd49f7c1",
   118 => x"86c487df",
   119 => x"c005a8c1",
   120 => x"d4ff87ea",
   121 => x"78ffc348",
   122 => x"c0c0c0c1",
   123 => x"c01ec0c0",
   124 => x"e9c1f0e1",
   125 => x"87c1fd49",
   126 => x"987086c4",
   127 => x"ff87ca05",
   128 => x"ffc348d4",
   129 => x"cb48c178",
   130 => x"87e6fe87",
   131 => x"fe058bc1",
   132 => x"48c087fd",
   133 => x"1e87defc",
   134 => x"d4ff1e73",
   135 => x"78ffc348",
   136 => x"1ec04bd3",
   137 => x"c1f0ffc0",
   138 => x"ccfc49c1",
   139 => x"7086c487",
   140 => x"87ca0598",
   141 => x"c348d4ff",
   142 => x"48c178ff",
   143 => x"f1fd87cb",
   144 => x"058bc187",
   145 => x"c087dbff",
   146 => x"87e9fb48",
   147 => x"5c5b5e0e",
   148 => x"4cd4ff0e",
   149 => x"c687dbfd",
   150 => x"e1c01eea",
   151 => x"49c8c1f0",
   152 => x"c487d6fb",
   153 => x"02a8c186",
   154 => x"eafe87c8",
   155 => x"c148c087",
   156 => x"d2fa87e2",
   157 => x"cf497087",
   158 => x"c699ffff",
   159 => x"c802a9ea",
   160 => x"87d3fe87",
   161 => x"cbc148c0",
   162 => x"7cffc387",
   163 => x"fc4bf1c0",
   164 => x"987087f4",
   165 => x"87ebc002",
   166 => x"ffc01ec0",
   167 => x"49fac1f0",
   168 => x"c487d6fa",
   169 => x"05987086",
   170 => x"ffc387d9",
   171 => x"c3496c7c",
   172 => x"7c7c7cff",
   173 => x"99c0c17c",
   174 => x"c187c402",
   175 => x"c087d548",
   176 => x"c287d148",
   177 => x"87c405ab",
   178 => x"87c848c0",
   179 => x"fe058bc1",
   180 => x"48c087fd",
   181 => x"1e87dcf9",
   182 => x"dbc21e73",
   183 => x"78c148cc",
   184 => x"d0ff4bc7",
   185 => x"fb78c248",
   186 => x"d0ff87c8",
   187 => x"c078c348",
   188 => x"d0e5c01e",
   189 => x"f849c0c1",
   190 => x"86c487ff",
   191 => x"c105a8c1",
   192 => x"abc24b87",
   193 => x"c087c505",
   194 => x"87f9c048",
   195 => x"ff058bc1",
   196 => x"f7fc87d0",
   197 => x"d0dbc287",
   198 => x"05987058",
   199 => x"1ec187cd",
   200 => x"c1f0ffc0",
   201 => x"d0f849d0",
   202 => x"ff86c487",
   203 => x"ffc348d4",
   204 => x"87ddc478",
   205 => x"58d4dbc2",
   206 => x"c248d0ff",
   207 => x"48d4ff78",
   208 => x"c178ffc3",
   209 => x"87edf748",
   210 => x"5c5b5e0e",
   211 => x"4a710e5d",
   212 => x"ff4dffc3",
   213 => x"7c754cd4",
   214 => x"c448d0ff",
   215 => x"7c7578c3",
   216 => x"ffc01e72",
   217 => x"49d8c1f0",
   218 => x"c487cef7",
   219 => x"02987086",
   220 => x"48c187c5",
   221 => x"7587eec0",
   222 => x"7cfec37c",
   223 => x"d41ec0c8",
   224 => x"f2f44966",
   225 => x"7586c487",
   226 => x"757c757c",
   227 => x"e0dad87c",
   228 => x"6c7c754b",
   229 => x"c187c505",
   230 => x"87f5058b",
   231 => x"d0ff7c75",
   232 => x"c078c248",
   233 => x"87c9f648",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"eec54cc0",
   237 => x"ff4adfcd",
   238 => x"ffc348d4",
   239 => x"c3486878",
   240 => x"c005a8fe",
   241 => x"d4ff87fe",
   242 => x"029b734d",
   243 => x"66d087cc",
   244 => x"f449731e",
   245 => x"86c487c8",
   246 => x"d0ff87d6",
   247 => x"78d1c448",
   248 => x"d07dffc3",
   249 => x"88c14866",
   250 => x"7058a6d4",
   251 => x"87f00598",
   252 => x"c348d4ff",
   253 => x"737878ff",
   254 => x"87c5059b",
   255 => x"d048d0ff",
   256 => x"4c4ac178",
   257 => x"fe058ac1",
   258 => x"487487ed",
   259 => x"1e87e2f4",
   260 => x"4a711e73",
   261 => x"d4ff4bc0",
   262 => x"78ffc348",
   263 => x"c448d0ff",
   264 => x"d4ff78c3",
   265 => x"78ffc348",
   266 => x"ffc01e72",
   267 => x"49d1c1f0",
   268 => x"c487c6f4",
   269 => x"05987086",
   270 => x"c0c887d2",
   271 => x"4966cc1e",
   272 => x"c487e5fd",
   273 => x"ff4b7086",
   274 => x"78c248d0",
   275 => x"e4f34873",
   276 => x"5b5e0e87",
   277 => x"c00e5d5c",
   278 => x"f0ffc01e",
   279 => x"f349c9c1",
   280 => x"1ed287d7",
   281 => x"49d4dbc2",
   282 => x"c887fdfc",
   283 => x"c14cc086",
   284 => x"acb7d284",
   285 => x"c287f804",
   286 => x"bf97d4db",
   287 => x"99c0c349",
   288 => x"05a9c0c1",
   289 => x"c287e7c0",
   290 => x"bf97dbdb",
   291 => x"c231d049",
   292 => x"bf97dcdb",
   293 => x"7232c84a",
   294 => x"dddbc2b1",
   295 => x"b14abf97",
   296 => x"ffcf4c71",
   297 => x"c19cffff",
   298 => x"c134ca84",
   299 => x"dbc287e7",
   300 => x"49bf97dd",
   301 => x"99c631c1",
   302 => x"97dedbc2",
   303 => x"b7c74abf",
   304 => x"c2b1722a",
   305 => x"bf97d9db",
   306 => x"9dcf4d4a",
   307 => x"97dadbc2",
   308 => x"9ac34abf",
   309 => x"dbc232ca",
   310 => x"4bbf97db",
   311 => x"b27333c2",
   312 => x"97dcdbc2",
   313 => x"c0c34bbf",
   314 => x"2bb7c69b",
   315 => x"81c2b273",
   316 => x"307148c1",
   317 => x"48c14970",
   318 => x"4d703075",
   319 => x"84c14c72",
   320 => x"c0c89471",
   321 => x"cc06adb7",
   322 => x"b734c187",
   323 => x"b7c0c82d",
   324 => x"f4ff01ad",
   325 => x"f0487487",
   326 => x"5e0e87d7",
   327 => x"0e5d5c5b",
   328 => x"e3c286f8",
   329 => x"78c048fa",
   330 => x"1ef2dbc2",
   331 => x"defb49c0",
   332 => x"7086c487",
   333 => x"87c50598",
   334 => x"c0c948c0",
   335 => x"c14dc087",
   336 => x"ddf2c07e",
   337 => x"dcc249bf",
   338 => x"c8714ae8",
   339 => x"87d9ec4b",
   340 => x"c2059870",
   341 => x"c07ec087",
   342 => x"49bfd9f2",
   343 => x"4ac4ddc2",
   344 => x"ec4bc871",
   345 => x"987087c3",
   346 => x"c087c205",
   347 => x"c0026e7e",
   348 => x"e2c287fd",
   349 => x"c24dbff8",
   350 => x"bf9ff0e3",
   351 => x"d6c5487e",
   352 => x"c705a8ea",
   353 => x"f8e2c287",
   354 => x"87ce4dbf",
   355 => x"e9ca486e",
   356 => x"c502a8d5",
   357 => x"c748c087",
   358 => x"dbc287e3",
   359 => x"49751ef2",
   360 => x"c487ecf9",
   361 => x"05987086",
   362 => x"48c087c5",
   363 => x"c087cec7",
   364 => x"49bfd9f2",
   365 => x"4ac4ddc2",
   366 => x"ea4bc871",
   367 => x"987087eb",
   368 => x"c287c805",
   369 => x"c148fae3",
   370 => x"c087da78",
   371 => x"49bfddf2",
   372 => x"4ae8dcc2",
   373 => x"ea4bc871",
   374 => x"987087cf",
   375 => x"87c5c002",
   376 => x"d8c648c0",
   377 => x"f0e3c287",
   378 => x"c149bf97",
   379 => x"c005a9d5",
   380 => x"e3c287cd",
   381 => x"49bf97f1",
   382 => x"02a9eac2",
   383 => x"c087c5c0",
   384 => x"87f9c548",
   385 => x"97f2dbc2",
   386 => x"c3487ebf",
   387 => x"c002a8e9",
   388 => x"486e87ce",
   389 => x"02a8ebc3",
   390 => x"c087c5c0",
   391 => x"87ddc548",
   392 => x"97fddbc2",
   393 => x"059949bf",
   394 => x"c287ccc0",
   395 => x"bf97fedb",
   396 => x"02a9c249",
   397 => x"c087c5c0",
   398 => x"87c1c548",
   399 => x"97ffdbc2",
   400 => x"e3c248bf",
   401 => x"4c7058f6",
   402 => x"c288c148",
   403 => x"c258fae3",
   404 => x"bf97c0dc",
   405 => x"c2817549",
   406 => x"bf97c1dc",
   407 => x"7232c84a",
   408 => x"e8c27ea1",
   409 => x"786e48c7",
   410 => x"97c2dcc2",
   411 => x"a6c848bf",
   412 => x"fae3c258",
   413 => x"cfc202bf",
   414 => x"d9f2c087",
   415 => x"ddc249bf",
   416 => x"c8714ac4",
   417 => x"87e1e74b",
   418 => x"c0029870",
   419 => x"48c087c5",
   420 => x"c287eac3",
   421 => x"4cbff2e3",
   422 => x"5cdbe8c2",
   423 => x"97d7dcc2",
   424 => x"31c849bf",
   425 => x"97d6dcc2",
   426 => x"49a14abf",
   427 => x"97d8dcc2",
   428 => x"32d04abf",
   429 => x"c249a172",
   430 => x"bf97d9dc",
   431 => x"7232d84a",
   432 => x"66c449a1",
   433 => x"c7e8c291",
   434 => x"e8c281bf",
   435 => x"dcc259cf",
   436 => x"4abf97df",
   437 => x"dcc232c8",
   438 => x"4bbf97de",
   439 => x"dcc24aa2",
   440 => x"4bbf97e0",
   441 => x"a27333d0",
   442 => x"e1dcc24a",
   443 => x"cf4bbf97",
   444 => x"7333d89b",
   445 => x"e8c24aa2",
   446 => x"8ac25ad3",
   447 => x"e8c29274",
   448 => x"a17248d3",
   449 => x"87c1c178",
   450 => x"97c4dcc2",
   451 => x"31c849bf",
   452 => x"97c3dcc2",
   453 => x"49a14abf",
   454 => x"ffc731c5",
   455 => x"c229c981",
   456 => x"c259dbe8",
   457 => x"bf97c9dc",
   458 => x"c232c84a",
   459 => x"bf97c8dc",
   460 => x"c44aa24b",
   461 => x"826e9266",
   462 => x"5ad7e8c2",
   463 => x"48cfe8c2",
   464 => x"e8c278c0",
   465 => x"a17248cb",
   466 => x"dbe8c278",
   467 => x"cfe8c248",
   468 => x"e8c278bf",
   469 => x"e8c248df",
   470 => x"c278bfd3",
   471 => x"02bffae3",
   472 => x"7487c9c0",
   473 => x"7030c448",
   474 => x"87c9c07e",
   475 => x"bfd7e8c2",
   476 => x"7030c448",
   477 => x"fee3c27e",
   478 => x"c1786e48",
   479 => x"268ef848",
   480 => x"264c264d",
   481 => x"0e4f264b",
   482 => x"5d5c5b5e",
   483 => x"c24a710e",
   484 => x"02bffae3",
   485 => x"4b7287cb",
   486 => x"4d722bc7",
   487 => x"c99dffc1",
   488 => x"c84b7287",
   489 => x"c34d722b",
   490 => x"e8c29dff",
   491 => x"c083bfc7",
   492 => x"abbfd5f2",
   493 => x"c087d902",
   494 => x"c25bd9f2",
   495 => x"731ef2db",
   496 => x"87cbf149",
   497 => x"987086c4",
   498 => x"c087c505",
   499 => x"87e6c048",
   500 => x"bffae3c2",
   501 => x"7587d202",
   502 => x"c291c449",
   503 => x"6981f2db",
   504 => x"ffffcf4c",
   505 => x"cb9cffff",
   506 => x"c2497587",
   507 => x"f2dbc291",
   508 => x"4c699f81",
   509 => x"c6fe4874",
   510 => x"5b5e0e87",
   511 => x"f80e5d5c",
   512 => x"9c4c7186",
   513 => x"c087c505",
   514 => x"87c0c348",
   515 => x"487ea4c8",
   516 => x"66d878c0",
   517 => x"d887c702",
   518 => x"05bf9766",
   519 => x"48c087c5",
   520 => x"c087e9c2",
   521 => x"4949c11e",
   522 => x"c487d3ca",
   523 => x"9d4d7086",
   524 => x"87c2c102",
   525 => x"4ac2e4c2",
   526 => x"e04966d8",
   527 => x"987087d0",
   528 => x"87f2c002",
   529 => x"66d84a75",
   530 => x"e04bcb49",
   531 => x"987087f5",
   532 => x"87e2c002",
   533 => x"9d751ec0",
   534 => x"c887c702",
   535 => x"78c048a6",
   536 => x"a6c887c5",
   537 => x"c878c148",
   538 => x"d1c94966",
   539 => x"7086c487",
   540 => x"fe059d4d",
   541 => x"9d7587fe",
   542 => x"87cec102",
   543 => x"6e49a5dc",
   544 => x"da786948",
   545 => x"a6c449a5",
   546 => x"78a4c448",
   547 => x"c448699f",
   548 => x"c2780866",
   549 => x"02bffae3",
   550 => x"a5d487d2",
   551 => x"49699f49",
   552 => x"99ffffc0",
   553 => x"30d04871",
   554 => x"87c27e70",
   555 => x"486e7ec0",
   556 => x"80bf66c4",
   557 => x"780866c4",
   558 => x"a4cc7cc0",
   559 => x"bf66c449",
   560 => x"49a4d079",
   561 => x"48c179c0",
   562 => x"48c087c2",
   563 => x"eefa8ef8",
   564 => x"5b5e0e87",
   565 => x"4c710e5c",
   566 => x"cbc1029c",
   567 => x"49a4c887",
   568 => x"c3c10269",
   569 => x"cc496c87",
   570 => x"80714866",
   571 => x"7058a6d0",
   572 => x"f6e3c2b9",
   573 => x"baff4abf",
   574 => x"99719972",
   575 => x"87e5c002",
   576 => x"6b4ba4c4",
   577 => x"87fff949",
   578 => x"e3c27b70",
   579 => x"6c49bff2",
   580 => x"cc7c7181",
   581 => x"e3c2b966",
   582 => x"ff4abff6",
   583 => x"719972ba",
   584 => x"dbff0599",
   585 => x"7c66cc87",
   586 => x"1e87d6f9",
   587 => x"4b711e73",
   588 => x"87c7029b",
   589 => x"6949a3c8",
   590 => x"c087c505",
   591 => x"87f6c048",
   592 => x"bfcbe8c2",
   593 => x"4aa3c449",
   594 => x"8ac24a6a",
   595 => x"bff2e3c2",
   596 => x"49a17292",
   597 => x"bff6e3c2",
   598 => x"729a6b4a",
   599 => x"f2c049a1",
   600 => x"66c859d9",
   601 => x"e6ea711e",
   602 => x"7086c487",
   603 => x"87c40598",
   604 => x"87c248c0",
   605 => x"caf848c1",
   606 => x"1e731e87",
   607 => x"029b4b71",
   608 => x"a3c887c7",
   609 => x"c5056949",
   610 => x"c048c087",
   611 => x"e8c287f6",
   612 => x"c449bfcb",
   613 => x"4a6a4aa3",
   614 => x"e3c28ac2",
   615 => x"7292bff2",
   616 => x"e3c249a1",
   617 => x"6b4abff6",
   618 => x"49a1729a",
   619 => x"59d9f2c0",
   620 => x"711e66c8",
   621 => x"c487d1e6",
   622 => x"05987086",
   623 => x"48c087c4",
   624 => x"48c187c2",
   625 => x"0e87fcf6",
   626 => x"5d5c5b5e",
   627 => x"4b711e0e",
   628 => x"734d66d4",
   629 => x"ccc1029b",
   630 => x"49a3c887",
   631 => x"c4c10269",
   632 => x"4ca3d087",
   633 => x"bff6e3c2",
   634 => x"6cb9ff49",
   635 => x"d47e994a",
   636 => x"cd06a966",
   637 => x"7c7bc087",
   638 => x"c44aa3cc",
   639 => x"796a49a3",
   640 => x"497287ca",
   641 => x"d499c0f8",
   642 => x"8d714d66",
   643 => x"29c94975",
   644 => x"49731e71",
   645 => x"c287fafa",
   646 => x"731ef2db",
   647 => x"87cbfc49",
   648 => x"66d486c8",
   649 => x"d6f5267c",
   650 => x"1e731e87",
   651 => x"029b4b71",
   652 => x"c287e4c0",
   653 => x"735bdfe8",
   654 => x"c28ac24a",
   655 => x"49bff2e3",
   656 => x"cbe8c292",
   657 => x"807248bf",
   658 => x"58e3e8c2",
   659 => x"30c44871",
   660 => x"58c2e4c2",
   661 => x"c287edc0",
   662 => x"c248dbe8",
   663 => x"78bfcfe8",
   664 => x"48dfe8c2",
   665 => x"bfd3e8c2",
   666 => x"fae3c278",
   667 => x"87c902bf",
   668 => x"bff2e3c2",
   669 => x"c731c449",
   670 => x"d7e8c287",
   671 => x"31c449bf",
   672 => x"59c2e4c2",
   673 => x"0e87fcf3",
   674 => x"0e5c5b5e",
   675 => x"4bc04a71",
   676 => x"c0029a72",
   677 => x"a2da87e0",
   678 => x"4b699f49",
   679 => x"bffae3c2",
   680 => x"d487cf02",
   681 => x"699f49a2",
   682 => x"ffc04c49",
   683 => x"34d09cff",
   684 => x"4cc087c2",
   685 => x"4973b374",
   686 => x"f387eefd",
   687 => x"5e0e87c3",
   688 => x"0e5d5c5b",
   689 => x"4a7186f4",
   690 => x"9a727ec0",
   691 => x"c287d802",
   692 => x"c048eedb",
   693 => x"e6dbc278",
   694 => x"dfe8c248",
   695 => x"dbc278bf",
   696 => x"e8c248ea",
   697 => x"c278bfdb",
   698 => x"c048cfe4",
   699 => x"fee3c250",
   700 => x"dbc249bf",
   701 => x"714abfee",
   702 => x"c9c403aa",
   703 => x"cf497287",
   704 => x"e9c00599",
   705 => x"d5f2c087",
   706 => x"e6dbc248",
   707 => x"dbc278bf",
   708 => x"dbc21ef2",
   709 => x"c249bfe6",
   710 => x"c148e6db",
   711 => x"e37178a1",
   712 => x"86c487ed",
   713 => x"48d1f2c0",
   714 => x"78f2dbc2",
   715 => x"f2c087cc",
   716 => x"c048bfd1",
   717 => x"f2c080e0",
   718 => x"dbc258d5",
   719 => x"c148bfee",
   720 => x"f2dbc280",
   721 => x"0c912758",
   722 => x"97bf0000",
   723 => x"029d4dbf",
   724 => x"c387e3c2",
   725 => x"c202ade5",
   726 => x"f2c087dc",
   727 => x"cb4bbfd1",
   728 => x"4c1149a3",
   729 => x"c105accf",
   730 => x"497587d2",
   731 => x"89c199df",
   732 => x"e4c291cd",
   733 => x"a3c181c2",
   734 => x"c351124a",
   735 => x"51124aa3",
   736 => x"124aa3c5",
   737 => x"4aa3c751",
   738 => x"a3c95112",
   739 => x"ce51124a",
   740 => x"51124aa3",
   741 => x"124aa3d0",
   742 => x"4aa3d251",
   743 => x"a3d45112",
   744 => x"d651124a",
   745 => x"51124aa3",
   746 => x"124aa3d8",
   747 => x"4aa3dc51",
   748 => x"a3de5112",
   749 => x"c151124a",
   750 => x"87fac07e",
   751 => x"99c84974",
   752 => x"87ebc005",
   753 => x"99d04974",
   754 => x"dc87d105",
   755 => x"cbc00266",
   756 => x"dc497387",
   757 => x"98700f66",
   758 => x"87d3c002",
   759 => x"c6c0056e",
   760 => x"c2e4c287",
   761 => x"c050c048",
   762 => x"48bfd1f2",
   763 => x"c287ddc2",
   764 => x"c048cfe4",
   765 => x"e3c27e50",
   766 => x"c249bffe",
   767 => x"4abfeedb",
   768 => x"fb04aa71",
   769 => x"e8c287f7",
   770 => x"c005bfdf",
   771 => x"e3c287c8",
   772 => x"c102bffa",
   773 => x"dbc287f4",
   774 => x"ed49bfea",
   775 => x"dbc287e9",
   776 => x"a6c458ee",
   777 => x"eadbc248",
   778 => x"e3c278bf",
   779 => x"c002bffa",
   780 => x"66c487d8",
   781 => x"ffffcf49",
   782 => x"a999f8ff",
   783 => x"87c5c002",
   784 => x"e1c04cc0",
   785 => x"c04cc187",
   786 => x"66c487dc",
   787 => x"f8ffcf49",
   788 => x"c002a999",
   789 => x"a6c887c8",
   790 => x"c078c048",
   791 => x"a6c887c5",
   792 => x"c878c148",
   793 => x"9c744c66",
   794 => x"87dec005",
   795 => x"c24966c4",
   796 => x"f2e3c289",
   797 => x"e8c291bf",
   798 => x"7148bfcb",
   799 => x"eadbc280",
   800 => x"eedbc258",
   801 => x"f978c048",
   802 => x"48c087e3",
   803 => x"eeeb8ef4",
   804 => x"00000087",
   805 => x"ffffff00",
   806 => x"000ca1ff",
   807 => x"000caa00",
   808 => x"54414600",
   809 => x"20203233",
   810 => x"41460020",
   811 => x"20363154",
   812 => x"1e002020",
   813 => x"c348d4ff",
   814 => x"486878ff",
   815 => x"ff1e4f26",
   816 => x"ffc348d4",
   817 => x"48d0ff78",
   818 => x"ff78e1c0",
   819 => x"78d448d4",
   820 => x"48e3e8c2",
   821 => x"50bfd4ff",
   822 => x"ff1e4f26",
   823 => x"e0c048d0",
   824 => x"1e4f2678",
   825 => x"7087ccff",
   826 => x"c6029949",
   827 => x"a9fbc087",
   828 => x"7187f105",
   829 => x"0e4f2648",
   830 => x"0e5c5b5e",
   831 => x"4cc04b71",
   832 => x"7087f0fe",
   833 => x"c0029949",
   834 => x"ecc087f9",
   835 => x"f2c002a9",
   836 => x"a9fbc087",
   837 => x"87ebc002",
   838 => x"acb766cc",
   839 => x"d087c703",
   840 => x"87c20266",
   841 => x"99715371",
   842 => x"c187c202",
   843 => x"87c3fe84",
   844 => x"02994970",
   845 => x"ecc087cd",
   846 => x"87c702a9",
   847 => x"05a9fbc0",
   848 => x"d087d5ff",
   849 => x"87c30266",
   850 => x"c07b97c0",
   851 => x"c405a9ec",
   852 => x"c54a7487",
   853 => x"c04a7487",
   854 => x"48728a0a",
   855 => x"4d2687c2",
   856 => x"4b264c26",
   857 => x"fd1e4f26",
   858 => x"497087c9",
   859 => x"aaf0c04a",
   860 => x"c087c904",
   861 => x"c301aaf9",
   862 => x"8af0c087",
   863 => x"04aac1c1",
   864 => x"dac187c9",
   865 => x"87c301aa",
   866 => x"728af7c0",
   867 => x"0e4f2648",
   868 => x"5d5c5b5e",
   869 => x"7186f80e",
   870 => x"fc4dc04c",
   871 => x"4bc087e0",
   872 => x"97eef8c0",
   873 => x"a9c049bf",
   874 => x"fc87cf04",
   875 => x"83c187f5",
   876 => x"97eef8c0",
   877 => x"06ab49bf",
   878 => x"f8c087f1",
   879 => x"02bf97ee",
   880 => x"eefb87cf",
   881 => x"99497087",
   882 => x"c087c602",
   883 => x"f105a9ec",
   884 => x"fb4bc087",
   885 => x"7e7087dd",
   886 => x"c887d8fb",
   887 => x"d2fb58a6",
   888 => x"c14a7087",
   889 => x"49a4c883",
   890 => x"6e496997",
   891 => x"87da05a9",
   892 => x"9749a4c9",
   893 => x"66c44969",
   894 => x"87ce05a9",
   895 => x"9749a4ca",
   896 => x"05aa4969",
   897 => x"4dc187c4",
   898 => x"486e87d4",
   899 => x"02a8ecc0",
   900 => x"486e87c8",
   901 => x"05a8fbc0",
   902 => x"4bc087c4",
   903 => x"9d754dc1",
   904 => x"87effe02",
   905 => x"7387f3fa",
   906 => x"fc8ef848",
   907 => x"0e0087f0",
   908 => x"5d5c5b5e",
   909 => x"7186f80e",
   910 => x"4bd4ff7e",
   911 => x"e8c21e6e",
   912 => x"f4e649e8",
   913 => x"7086c487",
   914 => x"eac40298",
   915 => x"d5e3c187",
   916 => x"496e4dbf",
   917 => x"c887f8fc",
   918 => x"987058a6",
   919 => x"c487c505",
   920 => x"78c148a6",
   921 => x"c548d0ff",
   922 => x"7bd5c178",
   923 => x"c14966c4",
   924 => x"c131c689",
   925 => x"bf97d3e3",
   926 => x"b071484a",
   927 => x"d0ff7b70",
   928 => x"c278c448",
   929 => x"bf97e3e8",
   930 => x"0299d049",
   931 => x"78c587d7",
   932 => x"c07bd6c1",
   933 => x"7bffc34a",
   934 => x"e0c082c1",
   935 => x"87f504aa",
   936 => x"c448d0ff",
   937 => x"7bffc378",
   938 => x"c548d0ff",
   939 => x"7bd3c178",
   940 => x"78c47bc1",
   941 => x"06adb7c0",
   942 => x"c287ebc2",
   943 => x"4cbff0e8",
   944 => x"c2029c8d",
   945 => x"dbc287c2",
   946 => x"a6c47ef2",
   947 => x"78c0c848",
   948 => x"acb7c08c",
   949 => x"c887c603",
   950 => x"c078a4c0",
   951 => x"e3e8c24c",
   952 => x"d049bf97",
   953 => x"87d00299",
   954 => x"e8c21ec0",
   955 => x"fae849e8",
   956 => x"7086c487",
   957 => x"87f5c04a",
   958 => x"1ef2dbc2",
   959 => x"49e8e8c2",
   960 => x"c487e8e8",
   961 => x"ff4a7086",
   962 => x"c5c848d0",
   963 => x"7bd4c178",
   964 => x"7bbf976e",
   965 => x"80c1486e",
   966 => x"66c47e70",
   967 => x"c888c148",
   968 => x"987058a6",
   969 => x"87e8ff05",
   970 => x"c448d0ff",
   971 => x"059a7278",
   972 => x"48c087c5",
   973 => x"c187c2c1",
   974 => x"e8e8c21e",
   975 => x"87d1e649",
   976 => x"9c7486c4",
   977 => x"87fefd05",
   978 => x"06adb7c0",
   979 => x"e8c287d1",
   980 => x"78c048e8",
   981 => x"78c080d0",
   982 => x"e8c280f4",
   983 => x"c078bff4",
   984 => x"fd01adb7",
   985 => x"d0ff87d5",
   986 => x"c178c548",
   987 => x"7bc07bd3",
   988 => x"48c178c4",
   989 => x"c087c2c0",
   990 => x"268ef848",
   991 => x"264c264d",
   992 => x"0e4f264b",
   993 => x"5d5c5b5e",
   994 => x"4b711e0e",
   995 => x"ab4d4cc0",
   996 => x"87e8c004",
   997 => x"1ecff6c0",
   998 => x"c4029d75",
   999 => x"c24ac087",
  1000 => x"724ac187",
  1001 => x"87d6ec49",
  1002 => x"7e7086c4",
  1003 => x"056e84c1",
  1004 => x"4c7387c2",
  1005 => x"ac7385c1",
  1006 => x"87d8ff06",
  1007 => x"fe26486e",
  1008 => x"5e0e87f9",
  1009 => x"710e5c5b",
  1010 => x"0266cc4b",
  1011 => x"c04c87d8",
  1012 => x"d8028cf0",
  1013 => x"c14a7487",
  1014 => x"87d1028a",
  1015 => x"87cd028a",
  1016 => x"87c9028a",
  1017 => x"497387d9",
  1018 => x"d287c4f9",
  1019 => x"c01e7487",
  1020 => x"d7d9c149",
  1021 => x"731e7487",
  1022 => x"cfd9c149",
  1023 => x"fd86c887",
  1024 => x"5e0e87fb",
  1025 => x"0e5d5c5b",
  1026 => x"494c711e",
  1027 => x"e9c291de",
  1028 => x"85714dd0",
  1029 => x"c1026d97",
  1030 => x"e8c287dc",
  1031 => x"7449bffc",
  1032 => x"defd7181",
  1033 => x"487e7087",
  1034 => x"f2c00298",
  1035 => x"c4e9c287",
  1036 => x"cb4a704b",
  1037 => x"eec1ff49",
  1038 => x"cb4b7487",
  1039 => x"e7e3c193",
  1040 => x"c183c483",
  1041 => x"747bfac1",
  1042 => x"efc1c149",
  1043 => x"c17b7587",
  1044 => x"bf97d4e3",
  1045 => x"e9c21e49",
  1046 => x"e5fd49c4",
  1047 => x"7486c487",
  1048 => x"d7c1c149",
  1049 => x"c149c087",
  1050 => x"c287f6c2",
  1051 => x"c048e4e8",
  1052 => x"de49c178",
  1053 => x"fc2687ca",
  1054 => x"6f4c87c1",
  1055 => x"6e696461",
  1056 => x"2e2e2e67",
  1057 => x"1e731e00",
  1058 => x"c2494a71",
  1059 => x"81bffce8",
  1060 => x"87effb71",
  1061 => x"029b4b70",
  1062 => x"e74987c4",
  1063 => x"e8c287e9",
  1064 => x"78c048fc",
  1065 => x"d7dd49c1",
  1066 => x"87d3fb87",
  1067 => x"c149c01e",
  1068 => x"2687eec1",
  1069 => x"4a711e4f",
  1070 => x"c191cb49",
  1071 => x"c881e7e3",
  1072 => x"c2481181",
  1073 => x"c258e8e8",
  1074 => x"c048fce8",
  1075 => x"dc49c178",
  1076 => x"4f2687ee",
  1077 => x"0299711e",
  1078 => x"e4c187d2",
  1079 => x"50c048fc",
  1080 => x"c2c180f7",
  1081 => x"e3c140f5",
  1082 => x"87ce78e0",
  1083 => x"48f8e4c1",
  1084 => x"78d9e3c1",
  1085 => x"c2c180fc",
  1086 => x"4f2678ec",
  1087 => x"5c5b5e0e",
  1088 => x"86f40e5d",
  1089 => x"4df2dbc2",
  1090 => x"a6c44cc0",
  1091 => x"c278c048",
  1092 => x"48bffce8",
  1093 => x"c106a8c0",
  1094 => x"dbc287c0",
  1095 => x"029848f2",
  1096 => x"c087f7c0",
  1097 => x"c81ecff6",
  1098 => x"87c70266",
  1099 => x"c048a6c4",
  1100 => x"c487c578",
  1101 => x"78c148a6",
  1102 => x"e64966c4",
  1103 => x"86c487c0",
  1104 => x"84c14d70",
  1105 => x"c14866c4",
  1106 => x"58a6c880",
  1107 => x"bffce8c2",
  1108 => x"87c603ac",
  1109 => x"ff059d75",
  1110 => x"4cc087c9",
  1111 => x"c3029d75",
  1112 => x"f6c087dc",
  1113 => x"66c81ecf",
  1114 => x"cc87c702",
  1115 => x"78c048a6",
  1116 => x"a6cc87c5",
  1117 => x"cc78c148",
  1118 => x"c1e54966",
  1119 => x"7086c487",
  1120 => x"0298487e",
  1121 => x"4987e4c2",
  1122 => x"699781cb",
  1123 => x"0299d049",
  1124 => x"7487d4c1",
  1125 => x"c191cb49",
  1126 => x"c181e7e3",
  1127 => x"c879c5c2",
  1128 => x"51ffc381",
  1129 => x"91de4974",
  1130 => x"4dd0e9c2",
  1131 => x"c1c28571",
  1132 => x"a5c17d97",
  1133 => x"51e0c049",
  1134 => x"97c2e4c2",
  1135 => x"87d202bf",
  1136 => x"a5c284c1",
  1137 => x"c2e4c24b",
  1138 => x"fe49db4a",
  1139 => x"c187d8fb",
  1140 => x"a5cd87d9",
  1141 => x"c151c049",
  1142 => x"4ba5c284",
  1143 => x"49cb4a6e",
  1144 => x"87c3fbfe",
  1145 => x"7487c4c1",
  1146 => x"c191cb49",
  1147 => x"c181e7e3",
  1148 => x"c279c2c0",
  1149 => x"bf97c2e4",
  1150 => x"7487d802",
  1151 => x"c191de49",
  1152 => x"d0e9c284",
  1153 => x"c283714b",
  1154 => x"dd4ac2e4",
  1155 => x"d6fafe49",
  1156 => x"7487d887",
  1157 => x"c293de4b",
  1158 => x"cb83d0e9",
  1159 => x"51c049a3",
  1160 => x"6e7384c1",
  1161 => x"fe49cb4a",
  1162 => x"c487fcf9",
  1163 => x"80c14866",
  1164 => x"c758a6c8",
  1165 => x"c5c003ac",
  1166 => x"fc056e87",
  1167 => x"487487e4",
  1168 => x"f6f48ef4",
  1169 => x"1e731e87",
  1170 => x"cb494b71",
  1171 => x"e7e3c191",
  1172 => x"4aa1c881",
  1173 => x"48d3e3c1",
  1174 => x"a1c95012",
  1175 => x"eef8c04a",
  1176 => x"ca501248",
  1177 => x"d4e3c181",
  1178 => x"c1501148",
  1179 => x"bf97d4e3",
  1180 => x"49c01e49",
  1181 => x"c287cbf5",
  1182 => x"de48e4e8",
  1183 => x"d549c178",
  1184 => x"f32687fe",
  1185 => x"5e0e87f9",
  1186 => x"0e5d5c5b",
  1187 => x"4d7186f4",
  1188 => x"c191cb49",
  1189 => x"c881e7e3",
  1190 => x"a1ca4aa1",
  1191 => x"48a6c47e",
  1192 => x"bfececc2",
  1193 => x"bf976e78",
  1194 => x"4c66c44b",
  1195 => x"48122c73",
  1196 => x"7058a6cc",
  1197 => x"c984c19c",
  1198 => x"49699781",
  1199 => x"c204acb7",
  1200 => x"6e4cc087",
  1201 => x"c84abf97",
  1202 => x"31724966",
  1203 => x"66c4b9ff",
  1204 => x"72487499",
  1205 => x"484a7030",
  1206 => x"ecc2b071",
  1207 => x"e5c058f0",
  1208 => x"49c087da",
  1209 => x"7587d9d4",
  1210 => x"cff7c049",
  1211 => x"f28ef487",
  1212 => x"731e87c9",
  1213 => x"494b711e",
  1214 => x"7387cbfe",
  1215 => x"87c6fe49",
  1216 => x"1e87fcf1",
  1217 => x"4b711e73",
  1218 => x"024aa3c6",
  1219 => x"c187e3c0",
  1220 => x"87d6028a",
  1221 => x"e8c1028a",
  1222 => x"c1028a87",
  1223 => x"028a87ca",
  1224 => x"8a87efc0",
  1225 => x"c187d902",
  1226 => x"49c787e9",
  1227 => x"c187c6f6",
  1228 => x"e8c287ec",
  1229 => x"78df48e4",
  1230 => x"c3d349c1",
  1231 => x"87dec187",
  1232 => x"bffce8c2",
  1233 => x"87cbc102",
  1234 => x"c288c148",
  1235 => x"c158c0e9",
  1236 => x"e9c287c1",
  1237 => x"c002bfc0",
  1238 => x"e8c287f9",
  1239 => x"c148bffc",
  1240 => x"c0e9c280",
  1241 => x"87ebc058",
  1242 => x"bffce8c2",
  1243 => x"c289c649",
  1244 => x"c059c0e9",
  1245 => x"da03a9b7",
  1246 => x"fce8c287",
  1247 => x"d278c048",
  1248 => x"c0e9c287",
  1249 => x"87cb02bf",
  1250 => x"bffce8c2",
  1251 => x"c280c648",
  1252 => x"c058c0e9",
  1253 => x"87e8d149",
  1254 => x"f4c04973",
  1255 => x"deef87de",
  1256 => x"5b5e0e87",
  1257 => x"ff0e5d5c",
  1258 => x"a6dc86d4",
  1259 => x"48a6c859",
  1260 => x"80c478c0",
  1261 => x"7866c0c1",
  1262 => x"78c180c4",
  1263 => x"78c180c4",
  1264 => x"48c0e9c2",
  1265 => x"e8c278c1",
  1266 => x"de48bfe4",
  1267 => x"87c905a8",
  1268 => x"cc87e9f4",
  1269 => x"e6cf58a6",
  1270 => x"87e2e387",
  1271 => x"e387c4e4",
  1272 => x"4c7087d1",
  1273 => x"02acfbc0",
  1274 => x"d887fbc1",
  1275 => x"edc10566",
  1276 => x"66fcc087",
  1277 => x"6a82c44a",
  1278 => x"c11e727e",
  1279 => x"c448f4df",
  1280 => x"a1c84966",
  1281 => x"7141204a",
  1282 => x"87f905aa",
  1283 => x"4a265110",
  1284 => x"4866fcc0",
  1285 => x"78c5c9c1",
  1286 => x"81c7496a",
  1287 => x"fcc05174",
  1288 => x"81c84966",
  1289 => x"fcc051c1",
  1290 => x"81c94966",
  1291 => x"fcc051c0",
  1292 => x"81ca4966",
  1293 => x"1ec151c0",
  1294 => x"496a1ed8",
  1295 => x"f6e281c8",
  1296 => x"c186c887",
  1297 => x"c04866c0",
  1298 => x"87c701a8",
  1299 => x"c148a6c8",
  1300 => x"c187ce78",
  1301 => x"c14866c0",
  1302 => x"58a6d088",
  1303 => x"c2e287c3",
  1304 => x"48a6d087",
  1305 => x"9c7478c2",
  1306 => x"87cfcd02",
  1307 => x"c14866c8",
  1308 => x"03a866c4",
  1309 => x"dc87c4cd",
  1310 => x"78c048a6",
  1311 => x"78c080e8",
  1312 => x"7087f0e0",
  1313 => x"acd0c14c",
  1314 => x"87d7c205",
  1315 => x"e37e66c4",
  1316 => x"a6c887d4",
  1317 => x"87dbe058",
  1318 => x"ecc04c70",
  1319 => x"edc105ac",
  1320 => x"4966c887",
  1321 => x"fcc091cb",
  1322 => x"a1c48166",
  1323 => x"c84d6a4a",
  1324 => x"66c44aa1",
  1325 => x"f5c2c152",
  1326 => x"f6dfff79",
  1327 => x"9c4c7087",
  1328 => x"c087d902",
  1329 => x"d302acfb",
  1330 => x"ff557487",
  1331 => x"7087e4df",
  1332 => x"c7029c4c",
  1333 => x"acfbc087",
  1334 => x"87edff05",
  1335 => x"c255e0c0",
  1336 => x"97c055c1",
  1337 => x"4866d87d",
  1338 => x"db05a86e",
  1339 => x"4866c887",
  1340 => x"04a866cc",
  1341 => x"66c887ca",
  1342 => x"cc80c148",
  1343 => x"87c858a6",
  1344 => x"c14866cc",
  1345 => x"58a6d088",
  1346 => x"87e7deff",
  1347 => x"d0c14c70",
  1348 => x"87c805ac",
  1349 => x"c14866d4",
  1350 => x"58a6d880",
  1351 => x"02acd0c1",
  1352 => x"c487e9fd",
  1353 => x"66d84866",
  1354 => x"e0c905a8",
  1355 => x"a6e0c087",
  1356 => x"7478c048",
  1357 => x"88fbc048",
  1358 => x"98487e70",
  1359 => x"87e2c902",
  1360 => x"7088cb48",
  1361 => x"0298487e",
  1362 => x"4887cdc1",
  1363 => x"7e7088c9",
  1364 => x"c3029848",
  1365 => x"c44887fe",
  1366 => x"487e7088",
  1367 => x"87ce0298",
  1368 => x"7088c148",
  1369 => x"0298487e",
  1370 => x"c887e9c3",
  1371 => x"a6dc87d6",
  1372 => x"78f0c048",
  1373 => x"87fbdcff",
  1374 => x"ecc04c70",
  1375 => x"c4c002ac",
  1376 => x"a6e0c087",
  1377 => x"acecc05c",
  1378 => x"ff87cd02",
  1379 => x"7087e4dc",
  1380 => x"acecc04c",
  1381 => x"87f3ff05",
  1382 => x"02acecc0",
  1383 => x"ff87c4c0",
  1384 => x"c087d0dc",
  1385 => x"d01eca1e",
  1386 => x"91cb4966",
  1387 => x"4866c4c1",
  1388 => x"a6cc8071",
  1389 => x"4866c858",
  1390 => x"a6d080c4",
  1391 => x"bf66cc58",
  1392 => x"f2dcff49",
  1393 => x"de1ec187",
  1394 => x"bf66d41e",
  1395 => x"e6dcff49",
  1396 => x"7086d087",
  1397 => x"08c04849",
  1398 => x"a6e8c088",
  1399 => x"06a8c058",
  1400 => x"c087eec0",
  1401 => x"dd4866e4",
  1402 => x"e4c003a8",
  1403 => x"bf66c487",
  1404 => x"66e4c049",
  1405 => x"51e0c081",
  1406 => x"4966e4c0",
  1407 => x"66c481c1",
  1408 => x"c1c281bf",
  1409 => x"66e4c051",
  1410 => x"c481c249",
  1411 => x"c081bf66",
  1412 => x"c1486e51",
  1413 => x"6e78c5c9",
  1414 => x"d081c849",
  1415 => x"496e5166",
  1416 => x"66d481c9",
  1417 => x"ca496e51",
  1418 => x"5166dc81",
  1419 => x"c14866d0",
  1420 => x"58a6d480",
  1421 => x"cc4866c8",
  1422 => x"c004a866",
  1423 => x"66c887cb",
  1424 => x"cc80c148",
  1425 => x"d9c558a6",
  1426 => x"4866cc87",
  1427 => x"a6d088c1",
  1428 => x"87cec558",
  1429 => x"87cedcff",
  1430 => x"58a6e8c0",
  1431 => x"87c6dcff",
  1432 => x"58a6e0c0",
  1433 => x"05a8ecc0",
  1434 => x"dc87cac0",
  1435 => x"e4c048a6",
  1436 => x"c4c07866",
  1437 => x"fad8ff87",
  1438 => x"4966c887",
  1439 => x"fcc091cb",
  1440 => x"80714866",
  1441 => x"c84a7e70",
  1442 => x"ca496e82",
  1443 => x"66e4c081",
  1444 => x"4966dc51",
  1445 => x"e4c081c1",
  1446 => x"48c18966",
  1447 => x"49703071",
  1448 => x"977189c1",
  1449 => x"ececc27a",
  1450 => x"e4c049bf",
  1451 => x"6a972966",
  1452 => x"9871484a",
  1453 => x"58a6ecc0",
  1454 => x"81c4496e",
  1455 => x"66d84d69",
  1456 => x"a866c448",
  1457 => x"87c8c002",
  1458 => x"c048a6c4",
  1459 => x"87c5c078",
  1460 => x"c148a6c4",
  1461 => x"1e66c478",
  1462 => x"751ee0c0",
  1463 => x"d6d8ff49",
  1464 => x"7086c887",
  1465 => x"acb7c04c",
  1466 => x"87d4c106",
  1467 => x"e0c08574",
  1468 => x"75897449",
  1469 => x"fddfc14b",
  1470 => x"e6fe714a",
  1471 => x"85c287e9",
  1472 => x"4866e0c0",
  1473 => x"e4c080c1",
  1474 => x"e8c058a6",
  1475 => x"81c14966",
  1476 => x"c002a970",
  1477 => x"a6c487c8",
  1478 => x"c078c048",
  1479 => x"a6c487c5",
  1480 => x"c478c148",
  1481 => x"a4c21e66",
  1482 => x"48e0c049",
  1483 => x"49708871",
  1484 => x"ff49751e",
  1485 => x"c887c0d7",
  1486 => x"a8b7c086",
  1487 => x"87c0ff01",
  1488 => x"0266e0c0",
  1489 => x"6e87d1c0",
  1490 => x"c081c949",
  1491 => x"6e5166e0",
  1492 => x"c6cac148",
  1493 => x"87ccc078",
  1494 => x"81c9496e",
  1495 => x"486e51c2",
  1496 => x"78f2cbc1",
  1497 => x"cc4866c8",
  1498 => x"c004a866",
  1499 => x"66c887cb",
  1500 => x"cc80c148",
  1501 => x"e9c058a6",
  1502 => x"4866cc87",
  1503 => x"a6d088c1",
  1504 => x"87dec058",
  1505 => x"87dbd5ff",
  1506 => x"d5c04c70",
  1507 => x"acc6c187",
  1508 => x"87c8c005",
  1509 => x"c14866d0",
  1510 => x"58a6d480",
  1511 => x"87c3d5ff",
  1512 => x"66d44c70",
  1513 => x"d880c148",
  1514 => x"9c7458a6",
  1515 => x"87cbc002",
  1516 => x"c14866c8",
  1517 => x"04a866c4",
  1518 => x"ff87fcf2",
  1519 => x"c887dbd4",
  1520 => x"a8c74866",
  1521 => x"87e5c003",
  1522 => x"48c0e9c2",
  1523 => x"66c878c0",
  1524 => x"c091cb49",
  1525 => x"c48166fc",
  1526 => x"4a6a4aa1",
  1527 => x"c87952c0",
  1528 => x"80c14866",
  1529 => x"c758a6cc",
  1530 => x"dbff04a8",
  1531 => x"8ed4ff87",
  1532 => x"87c7deff",
  1533 => x"64616f4c",
  1534 => x"202e2a20",
  1535 => x"00203a00",
  1536 => x"711e731e",
  1537 => x"c6029b4b",
  1538 => x"fce8c287",
  1539 => x"c778c048",
  1540 => x"fce8c21e",
  1541 => x"e3c11ebf",
  1542 => x"e8c21ee7",
  1543 => x"ed49bfe4",
  1544 => x"86cc87ff",
  1545 => x"bfe4e8c2",
  1546 => x"87e8e249",
  1547 => x"c8029b73",
  1548 => x"e7e3c187",
  1549 => x"d5e3c049",
  1550 => x"c2ddff87",
  1551 => x"e3c11e87",
  1552 => x"50c048d3",
  1553 => x"bfcae5c1",
  1554 => x"e2d7ff49",
  1555 => x"2648c087",
  1556 => x"d9c71e4f",
  1557 => x"fe49c187",
  1558 => x"e9c287e6",
  1559 => x"50c048c4",
  1560 => x"87f3e9fe",
  1561 => x"cd029870",
  1562 => x"edf2fe87",
  1563 => x"02987087",
  1564 => x"4ac187c4",
  1565 => x"4ac087c2",
  1566 => x"ce059a72",
  1567 => x"c11ec087",
  1568 => x"c049fde2",
  1569 => x"c487fbef",
  1570 => x"c287fe86",
  1571 => x"c048fce8",
  1572 => x"e4e8c278",
  1573 => x"1e78c048",
  1574 => x"49c8e3c1",
  1575 => x"87e2efc0",
  1576 => x"d8fe1ec0",
  1577 => x"c0497087",
  1578 => x"c887d7ef",
  1579 => x"87fdc286",
  1580 => x"87d7e3c0",
  1581 => x"87c4f3c0",
  1582 => x"2687f5ff",
  1583 => x"2044534f",
  1584 => x"6c696166",
  1585 => x"002e6465",
  1586 => x"746f6f42",
  1587 => x"2e676e69",
  1588 => x"00002e2e",
  1589 => x"00000100",
  1590 => x"45208000",
  1591 => x"00746978",
  1592 => x"61422080",
  1593 => x"02006b63",
  1594 => x"50000010",
  1595 => x"0000002a",
  1596 => x"10020000",
  1597 => x"2a6e0000",
  1598 => x"00000000",
  1599 => x"00100200",
  1600 => x"002a8c00",
  1601 => x"00000000",
  1602 => x"00001002",
  1603 => x"00002aaa",
  1604 => x"02000000",
  1605 => x"c8000010",
  1606 => x"0000002a",
  1607 => x"10020000",
  1608 => x"2ae60000",
  1609 => x"00000000",
  1610 => x"00100200",
  1611 => x"002b0400",
  1612 => x"00000000",
  1613 => x"000010b5",
  1614 => x"00000000",
  1615 => x"03000000",
  1616 => x"00000013",
  1617 => x"00000000",
  1618 => x"194e0000",
  1619 => x"4f420000",
  1620 => x"2020544f",
  1621 => x"4f522020",
  1622 => x"fe1e004d",
  1623 => x"78c048f0",
  1624 => x"097909cd",
  1625 => x"fe1e4f26",
  1626 => x"2648bff0",
  1627 => x"f0fe1e4f",
  1628 => x"2678c148",
  1629 => x"f0fe1e4f",
  1630 => x"2678c048",
  1631 => x"4a711e4f",
  1632 => x"265152c0",
  1633 => x"5b5e0e4f",
  1634 => x"f40e5d5c",
  1635 => x"974d7186",
  1636 => x"a5c17e6d",
  1637 => x"486c974c",
  1638 => x"6e58a6c8",
  1639 => x"a866c448",
  1640 => x"ff87c505",
  1641 => x"87e6c048",
  1642 => x"c287caff",
  1643 => x"6c9749a5",
  1644 => x"4ba3714b",
  1645 => x"974b6b97",
  1646 => x"486e7e6c",
  1647 => x"a6c880c1",
  1648 => x"cc98c758",
  1649 => x"977058a6",
  1650 => x"87e1fe7c",
  1651 => x"8ef44873",
  1652 => x"4c264d26",
  1653 => x"4f264b26",
  1654 => x"5c5b5e0e",
  1655 => x"7186f40e",
  1656 => x"4a66d84c",
  1657 => x"c29affc3",
  1658 => x"6c974ba4",
  1659 => x"49a17349",
  1660 => x"6c975172",
  1661 => x"c1486e7e",
  1662 => x"58a6c880",
  1663 => x"a6cc98c7",
  1664 => x"f4547058",
  1665 => x"87caff8e",
  1666 => x"e8fd1e1e",
  1667 => x"4abfe087",
  1668 => x"c0e0c049",
  1669 => x"87cb0299",
  1670 => x"ecc21e72",
  1671 => x"f7fe49e2",
  1672 => x"fd86c487",
  1673 => x"7e7087c0",
  1674 => x"2687c2fd",
  1675 => x"c21e4f26",
  1676 => x"fd49e2ec",
  1677 => x"e8c187c7",
  1678 => x"ddfc49c8",
  1679 => x"87eec387",
  1680 => x"5e0e4f26",
  1681 => x"0e5d5c5b",
  1682 => x"ecc24d71",
  1683 => x"f4fc49e2",
  1684 => x"c04b7087",
  1685 => x"c304abb7",
  1686 => x"f0c387c2",
  1687 => x"87c905ab",
  1688 => x"48e6ecc1",
  1689 => x"e3c278c1",
  1690 => x"abe0c387",
  1691 => x"c187c905",
  1692 => x"c148eaec",
  1693 => x"87d4c278",
  1694 => x"bfeaecc1",
  1695 => x"c287c602",
  1696 => x"c24ca3c0",
  1697 => x"c14c7387",
  1698 => x"02bfe6ec",
  1699 => x"7487e0c0",
  1700 => x"29b7c449",
  1701 => x"fdedc191",
  1702 => x"cf4a7481",
  1703 => x"c192c29a",
  1704 => x"70307248",
  1705 => x"72baff4a",
  1706 => x"70986948",
  1707 => x"7487db79",
  1708 => x"29b7c449",
  1709 => x"fdedc191",
  1710 => x"cf4a7481",
  1711 => x"c392c29a",
  1712 => x"70307248",
  1713 => x"b069484a",
  1714 => x"9d757970",
  1715 => x"87f0c005",
  1716 => x"c848d0ff",
  1717 => x"d4ff78e1",
  1718 => x"c178c548",
  1719 => x"02bfeaec",
  1720 => x"e0c387c3",
  1721 => x"e6ecc178",
  1722 => x"87c602bf",
  1723 => x"c348d4ff",
  1724 => x"d4ff78f0",
  1725 => x"ff0b7b0b",
  1726 => x"e1c848d0",
  1727 => x"78e0c078",
  1728 => x"48eaecc1",
  1729 => x"ecc178c0",
  1730 => x"78c048e6",
  1731 => x"49e2ecc2",
  1732 => x"7087f2f9",
  1733 => x"abb7c04b",
  1734 => x"87fefc03",
  1735 => x"4d2648c0",
  1736 => x"4b264c26",
  1737 => x"00004f26",
  1738 => x"00000000",
  1739 => x"c01e0000",
  1740 => x"c449724a",
  1741 => x"fdedc191",
  1742 => x"c179c081",
  1743 => x"aab7d082",
  1744 => x"2687ee04",
  1745 => x"5b5e0e4f",
  1746 => x"710e5d5c",
  1747 => x"87e5f84d",
  1748 => x"b7c44a75",
  1749 => x"edc1922a",
  1750 => x"4c7582fd",
  1751 => x"94c29ccf",
  1752 => x"744b496a",
  1753 => x"c29bc32b",
  1754 => x"70307448",
  1755 => x"74bcff4c",
  1756 => x"70987148",
  1757 => x"87f5f77a",
  1758 => x"e1fe4873",
  1759 => x"00000087",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"d0ff1e00",
  1776 => x"78e1c848",
  1777 => x"d4ff4871",
  1778 => x"4f267808",
  1779 => x"48d0ff1e",
  1780 => x"7178e1c8",
  1781 => x"08d4ff48",
  1782 => x"4866c478",
  1783 => x"7808d4ff",
  1784 => x"711e4f26",
  1785 => x"4966c44a",
  1786 => x"ff49721e",
  1787 => x"d0ff87de",
  1788 => x"78e0c048",
  1789 => x"1e4f2626",
  1790 => x"4b711e73",
  1791 => x"1e4966c8",
  1792 => x"e0c14a73",
  1793 => x"d9ff49a2",
  1794 => x"87c42687",
  1795 => x"4c264d26",
  1796 => x"4f264b26",
  1797 => x"711e731e",
  1798 => x"b7c24b4a",
  1799 => x"87c803ab",
  1800 => x"c34a49a3",
  1801 => x"87c79aff",
  1802 => x"4a49a3ce",
  1803 => x"c89affc3",
  1804 => x"721e4966",
  1805 => x"87eafe49",
  1806 => x"87d4ff26",
  1807 => x"4ad4ff1e",
  1808 => x"ff7affc3",
  1809 => x"e1c048d0",
  1810 => x"c27ade78",
  1811 => x"7abfecec",
  1812 => x"28c84849",
  1813 => x"48717a70",
  1814 => x"7a7028d0",
  1815 => x"28d84871",
  1816 => x"d0ff7a70",
  1817 => x"78e0c048",
  1818 => x"ff1e4f26",
  1819 => x"c9c848d0",
  1820 => x"ff487178",
  1821 => x"267808d4",
  1822 => x"4a711e4f",
  1823 => x"ff87eb49",
  1824 => x"78c848d0",
  1825 => x"731e4f26",
  1826 => x"c24b711e",
  1827 => x"02bffcec",
  1828 => x"ebc287c3",
  1829 => x"48d0ff87",
  1830 => x"7378c9c8",
  1831 => x"b0e0c048",
  1832 => x"7808d4ff",
  1833 => x"48f0ecc2",
  1834 => x"66c878c0",
  1835 => x"c387c502",
  1836 => x"87c249ff",
  1837 => x"ecc249c0",
  1838 => x"66cc59f8",
  1839 => x"c587c602",
  1840 => x"c44ad5d5",
  1841 => x"ffffcf87",
  1842 => x"fcecc24a",
  1843 => x"fcecc25a",
  1844 => x"c478c148",
  1845 => x"264d2687",
  1846 => x"264b264c",
  1847 => x"5b5e0e4f",
  1848 => x"710e5d5c",
  1849 => x"f8ecc24a",
  1850 => x"9a724cbf",
  1851 => x"4987cb02",
  1852 => x"f1c191c8",
  1853 => x"83714bfc",
  1854 => x"f5c187c4",
  1855 => x"4dc04bfc",
  1856 => x"99744913",
  1857 => x"bff4ecc2",
  1858 => x"ffb87148",
  1859 => x"c17808d4",
  1860 => x"c8852cb7",
  1861 => x"e704adb7",
  1862 => x"f0ecc287",
  1863 => x"80c848bf",
  1864 => x"58f4ecc2",
  1865 => x"1e87eefe",
  1866 => x"4b711e73",
  1867 => x"029a4a13",
  1868 => x"497287cb",
  1869 => x"1387e6fe",
  1870 => x"f5059a4a",
  1871 => x"87d9fe87",
  1872 => x"f0ecc21e",
  1873 => x"ecc249bf",
  1874 => x"a1c148f0",
  1875 => x"b7c0c478",
  1876 => x"87db03a9",
  1877 => x"c248d4ff",
  1878 => x"78bff4ec",
  1879 => x"bff0ecc2",
  1880 => x"f0ecc249",
  1881 => x"78a1c148",
  1882 => x"a9b7c0c4",
  1883 => x"ff87e504",
  1884 => x"78c848d0",
  1885 => x"48fcecc2",
  1886 => x"4f2678c0",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"5f000000",
  1890 => x"0000005f",
  1891 => x"00030300",
  1892 => x"00000303",
  1893 => x"147f7f14",
  1894 => x"00147f7f",
  1895 => x"6b2e2400",
  1896 => x"00123a6b",
  1897 => x"18366a4c",
  1898 => x"0032566c",
  1899 => x"594f7e30",
  1900 => x"40683a77",
  1901 => x"07040000",
  1902 => x"00000003",
  1903 => x"3e1c0000",
  1904 => x"00004163",
  1905 => x"63410000",
  1906 => x"00001c3e",
  1907 => x"1c3e2a08",
  1908 => x"082a3e1c",
  1909 => x"3e080800",
  1910 => x"0008083e",
  1911 => x"e0800000",
  1912 => x"00000060",
  1913 => x"08080800",
  1914 => x"00080808",
  1915 => x"60000000",
  1916 => x"00000060",
  1917 => x"18306040",
  1918 => x"0103060c",
  1919 => x"597f3e00",
  1920 => x"003e7f4d",
  1921 => x"7f060400",
  1922 => x"0000007f",
  1923 => x"71634200",
  1924 => x"00464f59",
  1925 => x"49632200",
  1926 => x"00367f49",
  1927 => x"13161c18",
  1928 => x"00107f7f",
  1929 => x"45672700",
  1930 => x"00397d45",
  1931 => x"4b7e3c00",
  1932 => x"00307949",
  1933 => x"71010100",
  1934 => x"00070f79",
  1935 => x"497f3600",
  1936 => x"00367f49",
  1937 => x"494f0600",
  1938 => x"001e3f69",
  1939 => x"66000000",
  1940 => x"00000066",
  1941 => x"e6800000",
  1942 => x"00000066",
  1943 => x"14080800",
  1944 => x"00222214",
  1945 => x"14141400",
  1946 => x"00141414",
  1947 => x"14222200",
  1948 => x"00080814",
  1949 => x"51030200",
  1950 => x"00060f59",
  1951 => x"5d417f3e",
  1952 => x"001e1f55",
  1953 => x"097f7e00",
  1954 => x"007e7f09",
  1955 => x"497f7f00",
  1956 => x"00367f49",
  1957 => x"633e1c00",
  1958 => x"00414141",
  1959 => x"417f7f00",
  1960 => x"001c3e63",
  1961 => x"497f7f00",
  1962 => x"00414149",
  1963 => x"097f7f00",
  1964 => x"00010109",
  1965 => x"417f3e00",
  1966 => x"007a7b49",
  1967 => x"087f7f00",
  1968 => x"007f7f08",
  1969 => x"7f410000",
  1970 => x"0000417f",
  1971 => x"40602000",
  1972 => x"003f7f40",
  1973 => x"1c087f7f",
  1974 => x"00416336",
  1975 => x"407f7f00",
  1976 => x"00404040",
  1977 => x"0c067f7f",
  1978 => x"007f7f06",
  1979 => x"0c067f7f",
  1980 => x"007f7f18",
  1981 => x"417f3e00",
  1982 => x"003e7f41",
  1983 => x"097f7f00",
  1984 => x"00060f09",
  1985 => x"61417f3e",
  1986 => x"00407e7f",
  1987 => x"097f7f00",
  1988 => x"00667f19",
  1989 => x"4d6f2600",
  1990 => x"00327b59",
  1991 => x"7f010100",
  1992 => x"0001017f",
  1993 => x"407f3f00",
  1994 => x"003f7f40",
  1995 => x"703f0f00",
  1996 => x"000f3f70",
  1997 => x"18307f7f",
  1998 => x"007f7f30",
  1999 => x"1c366341",
  2000 => x"4163361c",
  2001 => x"7c060301",
  2002 => x"0103067c",
  2003 => x"4d597161",
  2004 => x"00414347",
  2005 => x"7f7f0000",
  2006 => x"00004141",
  2007 => x"0c060301",
  2008 => x"40603018",
  2009 => x"41410000",
  2010 => x"00007f7f",
  2011 => x"03060c08",
  2012 => x"00080c06",
  2013 => x"80808080",
  2014 => x"00808080",
  2015 => x"03000000",
  2016 => x"00000407",
  2017 => x"54742000",
  2018 => x"00787c54",
  2019 => x"447f7f00",
  2020 => x"00387c44",
  2021 => x"447c3800",
  2022 => x"00004444",
  2023 => x"447c3800",
  2024 => x"007f7f44",
  2025 => x"547c3800",
  2026 => x"00185c54",
  2027 => x"7f7e0400",
  2028 => x"00000505",
  2029 => x"a4bc1800",
  2030 => x"007cfca4",
  2031 => x"047f7f00",
  2032 => x"00787c04",
  2033 => x"3d000000",
  2034 => x"0000407d",
  2035 => x"80808000",
  2036 => x"00007dfd",
  2037 => x"107f7f00",
  2038 => x"00446c38",
  2039 => x"3f000000",
  2040 => x"0000407f",
  2041 => x"180c7c7c",
  2042 => x"00787c0c",
  2043 => x"047c7c00",
  2044 => x"00787c04",
  2045 => x"447c3800",
  2046 => x"00387c44",
  2047 => x"24fcfc00",
  2048 => x"00183c24",
  2049 => x"243c1800",
  2050 => x"00fcfc24",
  2051 => x"047c7c00",
  2052 => x"00080c04",
  2053 => x"545c4800",
  2054 => x"00207454",
  2055 => x"7f3f0400",
  2056 => x"00004444",
  2057 => x"407c3c00",
  2058 => x"007c7c40",
  2059 => x"603c1c00",
  2060 => x"001c3c60",
  2061 => x"30607c3c",
  2062 => x"003c7c60",
  2063 => x"10386c44",
  2064 => x"00446c38",
  2065 => x"e0bc1c00",
  2066 => x"001c3c60",
  2067 => x"74644400",
  2068 => x"00444c5c",
  2069 => x"3e080800",
  2070 => x"00414177",
  2071 => x"7f000000",
  2072 => x"0000007f",
  2073 => x"77414100",
  2074 => x"0008083e",
  2075 => x"03010102",
  2076 => x"00010202",
  2077 => x"7f7f7f7f",
  2078 => x"007f7f7f",
  2079 => x"1c1c0808",
  2080 => x"7f7f3e3e",
  2081 => x"3e3e7f7f",
  2082 => x"08081c1c",
  2083 => x"7c181000",
  2084 => x"0010187c",
  2085 => x"7c301000",
  2086 => x"0010307c",
  2087 => x"60603010",
  2088 => x"00061e78",
  2089 => x"183c6642",
  2090 => x"0042663c",
  2091 => x"c26a3878",
  2092 => x"00386cc6",
  2093 => x"60000060",
  2094 => x"00600000",
  2095 => x"5c5b5e0e",
  2096 => x"711e0e5d",
  2097 => x"c1edc24c",
  2098 => x"4bc04dbf",
  2099 => x"ab741ec0",
  2100 => x"c487c702",
  2101 => x"78c048a6",
  2102 => x"a6c487c5",
  2103 => x"c478c148",
  2104 => x"49731e66",
  2105 => x"c887dfee",
  2106 => x"49e0c086",
  2107 => x"c487eeef",
  2108 => x"496a4aa5",
  2109 => x"f187f0f0",
  2110 => x"85cb87c6",
  2111 => x"b7c883c1",
  2112 => x"c7ff04ab",
  2113 => x"4d262687",
  2114 => x"4b264c26",
  2115 => x"711e4f26",
  2116 => x"c5edc24a",
  2117 => x"c5edc25a",
  2118 => x"4978c748",
  2119 => x"2687ddfe",
  2120 => x"1e731e4f",
  2121 => x"b7c04a71",
  2122 => x"87d303aa",
  2123 => x"bfdbd3c2",
  2124 => x"c187c405",
  2125 => x"c087c24b",
  2126 => x"dfd3c24b",
  2127 => x"c287c45b",
  2128 => x"c25adfd3",
  2129 => x"4abfdbd3",
  2130 => x"c0c19ac1",
  2131 => x"e8ec49a2",
  2132 => x"c248fc87",
  2133 => x"78bfdbd3",
  2134 => x"1e87effe",
  2135 => x"66c44a71",
  2136 => x"ea49721e",
  2137 => x"262687ee",
  2138 => x"d4ff1e4f",
  2139 => x"78ffc348",
  2140 => x"c048d0ff",
  2141 => x"d4ff78e1",
  2142 => x"7178c148",
  2143 => x"ff30c448",
  2144 => x"ff7808d4",
  2145 => x"e0c048d0",
  2146 => x"0e4f2678",
  2147 => x"5d5c5b5e",
  2148 => x"c486f40e",
  2149 => x"78c048a6",
  2150 => x"7ebfec4b",
  2151 => x"bfc1edc2",
  2152 => x"4cbfe84d",
  2153 => x"bfdbd3c2",
  2154 => x"87d6e249",
  2155 => x"cc49eecb",
  2156 => x"a6cc87f1",
  2157 => x"e649c758",
  2158 => x"987087cb",
  2159 => x"6e87c805",
  2160 => x"0299c149",
  2161 => x"c187c3c1",
  2162 => x"7ebfec4b",
  2163 => x"bfdbd3c2",
  2164 => x"87eee149",
  2165 => x"cc4966c8",
  2166 => x"987087d5",
  2167 => x"c287d802",
  2168 => x"49bfd3d3",
  2169 => x"d3c2b9c1",
  2170 => x"fd7159d7",
  2171 => x"eecb87fb",
  2172 => x"87efcb49",
  2173 => x"c758a6cc",
  2174 => x"87c9e549",
  2175 => x"ff059870",
  2176 => x"496e87c5",
  2177 => x"fe0599c1",
  2178 => x"9b7387fd",
  2179 => x"ff87d002",
  2180 => x"87cdfc49",
  2181 => x"e449dac1",
  2182 => x"a6c487eb",
  2183 => x"c278c148",
  2184 => x"05bfdbd3",
  2185 => x"c387e9c0",
  2186 => x"d8e449fd",
  2187 => x"49fac387",
  2188 => x"7487d2e4",
  2189 => x"99ffc349",
  2190 => x"49c01e71",
  2191 => x"7487dcfc",
  2192 => x"29b7c849",
  2193 => x"49c11e71",
  2194 => x"c887d0fc",
  2195 => x"87edc886",
  2196 => x"ffc34974",
  2197 => x"2cb7c899",
  2198 => x"9c74b471",
  2199 => x"c287dd02",
  2200 => x"49bfd7d3",
  2201 => x"7087c8ca",
  2202 => x"87c40598",
  2203 => x"87d24cc0",
  2204 => x"c949e0c2",
  2205 => x"d3c287ed",
  2206 => x"87c658db",
  2207 => x"48d7d3c2",
  2208 => x"497478c0",
  2209 => x"cd0599c2",
  2210 => x"49ebc387",
  2211 => x"7087f6e2",
  2212 => x"0299c249",
  2213 => x"d8c187cf",
  2214 => x"bf6e7ea5",
  2215 => x"87c5c002",
  2216 => x"7349fb4b",
  2217 => x"c149740f",
  2218 => x"87cd0599",
  2219 => x"e249f4c3",
  2220 => x"497087d3",
  2221 => x"cf0299c2",
  2222 => x"a5d8c187",
  2223 => x"02bf6e7e",
  2224 => x"4b87c5c0",
  2225 => x"0f7349fa",
  2226 => x"99c84974",
  2227 => x"c387ce05",
  2228 => x"f0e149f5",
  2229 => x"c2497087",
  2230 => x"e5c00299",
  2231 => x"c5edc287",
  2232 => x"cac002bf",
  2233 => x"88c14887",
  2234 => x"58c9edc2",
  2235 => x"c187cec0",
  2236 => x"6a4aa5d8",
  2237 => x"87c5c002",
  2238 => x"7349ff4b",
  2239 => x"48a6c40f",
  2240 => x"497478c1",
  2241 => x"c00599c4",
  2242 => x"f2c387ce",
  2243 => x"87f5e049",
  2244 => x"99c24970",
  2245 => x"87ecc002",
  2246 => x"bfc5edc2",
  2247 => x"b7c7487e",
  2248 => x"cbc003a8",
  2249 => x"c1486e87",
  2250 => x"c9edc280",
  2251 => x"87cfc058",
  2252 => x"7ea5d8c1",
  2253 => x"c002bf6e",
  2254 => x"fe4b87c5",
  2255 => x"c40f7349",
  2256 => x"78c148a6",
  2257 => x"ff49fdc3",
  2258 => x"7087fadf",
  2259 => x"0299c249",
  2260 => x"c287e5c0",
  2261 => x"02bfc5ed",
  2262 => x"c287c9c0",
  2263 => x"c048c5ed",
  2264 => x"87cfc078",
  2265 => x"7ea5d8c1",
  2266 => x"c002bf6e",
  2267 => x"fd4b87c5",
  2268 => x"c40f7349",
  2269 => x"78c148a6",
  2270 => x"ff49fac3",
  2271 => x"7087c6df",
  2272 => x"0299c249",
  2273 => x"c287e9c0",
  2274 => x"48bfc5ed",
  2275 => x"03a8b7c7",
  2276 => x"c287c9c0",
  2277 => x"c748c5ed",
  2278 => x"87cfc078",
  2279 => x"7ea5d8c1",
  2280 => x"c002bf6e",
  2281 => x"fc4b87c5",
  2282 => x"c40f7349",
  2283 => x"78c148a6",
  2284 => x"edc24bc0",
  2285 => x"50c048c0",
  2286 => x"c449eecb",
  2287 => x"a6cc87e5",
  2288 => x"c0edc258",
  2289 => x"c105bf97",
  2290 => x"497487de",
  2291 => x"0599f0c3",
  2292 => x"c187cdc0",
  2293 => x"ddff49da",
  2294 => x"987087eb",
  2295 => x"87c8c102",
  2296 => x"bfe84bc1",
  2297 => x"ffc3494c",
  2298 => x"2cb7c899",
  2299 => x"d3c2b471",
  2300 => x"ff49bfdb",
  2301 => x"c887cbd9",
  2302 => x"f2c34966",
  2303 => x"02987087",
  2304 => x"c287c6c0",
  2305 => x"c148c0ed",
  2306 => x"c0edc250",
  2307 => x"c005bf97",
  2308 => x"497487d6",
  2309 => x"0599f0c3",
  2310 => x"c187c5ff",
  2311 => x"dcff49da",
  2312 => x"987087e3",
  2313 => x"87f8fe05",
  2314 => x"c0029b73",
  2315 => x"a6c887dc",
  2316 => x"c5edc248",
  2317 => x"66c878bf",
  2318 => x"7591cb49",
  2319 => x"bf6e7ea1",
  2320 => x"87c6c002",
  2321 => x"4966c84b",
  2322 => x"66c40f73",
  2323 => x"87c8c002",
  2324 => x"bfc5edc2",
  2325 => x"87e4f149",
  2326 => x"bfdfd3c2",
  2327 => x"87ddc002",
  2328 => x"87cbc249",
  2329 => x"c0029870",
  2330 => x"edc287d3",
  2331 => x"f149bfc5",
  2332 => x"49c087ca",
  2333 => x"c287eaf2",
  2334 => x"c048dfd3",
  2335 => x"f28ef478",
  2336 => x"5e0e87c4",
  2337 => x"0e5d5c5b",
  2338 => x"c24c711e",
  2339 => x"49bfc1ed",
  2340 => x"4da1cdc1",
  2341 => x"6981d1c1",
  2342 => x"029c747e",
  2343 => x"a5c487cf",
  2344 => x"c27b744b",
  2345 => x"49bfc1ed",
  2346 => x"6e87e3f1",
  2347 => x"059c747b",
  2348 => x"4bc087c4",
  2349 => x"4bc187c2",
  2350 => x"e4f14973",
  2351 => x"0266d487",
  2352 => x"de4987c7",
  2353 => x"c24a7087",
  2354 => x"c24ac087",
  2355 => x"265ae3d3",
  2356 => x"0087f3f0",
  2357 => x"00000000",
  2358 => x"00000000",
  2359 => x"00000000",
  2360 => x"1e000000",
  2361 => x"c8ff4a71",
  2362 => x"a17249bf",
  2363 => x"1e4f2648",
  2364 => x"89bfc8ff",
  2365 => x"c0c0c0fe",
  2366 => x"01a9c0c0",
  2367 => x"4ac087c4",
  2368 => x"4ac187c2",
  2369 => x"4f264872",
  2370 => x"5c5b5e0e",
  2371 => x"4b710e5d",
  2372 => x"d04cd4ff",
  2373 => x"78c04866",
  2374 => x"daff49d6",
  2375 => x"ffc387df",
  2376 => x"c3496c7c",
  2377 => x"4d7199ff",
  2378 => x"99f0c349",
  2379 => x"05a9e0c1",
  2380 => x"ffc387cb",
  2381 => x"c3486c7c",
  2382 => x"0866d098",
  2383 => x"7cffc378",
  2384 => x"c8494a6c",
  2385 => x"7cffc331",
  2386 => x"b2714a6c",
  2387 => x"31c84972",
  2388 => x"6c7cffc3",
  2389 => x"72b2714a",
  2390 => x"c331c849",
  2391 => x"4a6c7cff",
  2392 => x"d0ffb271",
  2393 => x"78e0c048",
  2394 => x"c2029b73",
  2395 => x"757b7287",
  2396 => x"264d2648",
  2397 => x"264b264c",
  2398 => x"4f261e4f",
  2399 => x"5c5b5e0e",
  2400 => x"7686f80e",
  2401 => x"49a6c81e",
  2402 => x"c487fdfd",
  2403 => x"6e4b7086",
  2404 => x"01a8c048",
  2405 => x"7387f0c2",
  2406 => x"9af0c34a",
  2407 => x"02aad0c1",
  2408 => x"e0c187c7",
  2409 => x"dec205aa",
  2410 => x"c8497387",
  2411 => x"87c30299",
  2412 => x"7387c6ff",
  2413 => x"c29cc34c",
  2414 => x"c2c105ac",
  2415 => x"4966c487",
  2416 => x"1e7131c9",
  2417 => x"d44a66c4",
  2418 => x"c9edc292",
  2419 => x"fe817249",
  2420 => x"d887f4cf",
  2421 => x"e4d7ff49",
  2422 => x"1ec0c887",
  2423 => x"49f2dbc2",
  2424 => x"87faebfd",
  2425 => x"c048d0ff",
  2426 => x"dbc278e0",
  2427 => x"66cc1ef2",
  2428 => x"c292d44a",
  2429 => x"7249c9ed",
  2430 => x"fccdfe81",
  2431 => x"c186cc87",
  2432 => x"c2c105ac",
  2433 => x"4966c487",
  2434 => x"1e7131c9",
  2435 => x"d44a66c4",
  2436 => x"c9edc292",
  2437 => x"fe817249",
  2438 => x"c287ecce",
  2439 => x"c81ef2db",
  2440 => x"92d44a66",
  2441 => x"49c9edc2",
  2442 => x"cbfe8172",
  2443 => x"49d787fd",
  2444 => x"87c9d6ff",
  2445 => x"c21ec0c8",
  2446 => x"fd49f2db",
  2447 => x"cc87f8e9",
  2448 => x"48d0ff86",
  2449 => x"f878e0c0",
  2450 => x"87e7fc8e",
  2451 => x"5c5b5e0e",
  2452 => x"4a710e5d",
  2453 => x"d04cd4ff",
  2454 => x"b7c34d66",
  2455 => x"87c506ad",
  2456 => x"e1c148c0",
  2457 => x"751e7287",
  2458 => x"c293d44b",
  2459 => x"7383c9ed",
  2460 => x"c4c6fe49",
  2461 => x"6b83c887",
  2462 => x"48d0ff4b",
  2463 => x"dd78e1c8",
  2464 => x"c348737c",
  2465 => x"7c7098ff",
  2466 => x"b7c84973",
  2467 => x"c3487129",
  2468 => x"7c7098ff",
  2469 => x"b7d04973",
  2470 => x"c3487129",
  2471 => x"7c7098ff",
  2472 => x"b7d84873",
  2473 => x"c07c7028",
  2474 => x"7c7c7c7c",
  2475 => x"7c7c7c7c",
  2476 => x"7c7c7c7c",
  2477 => x"c048d0ff",
  2478 => x"1e7578e0",
  2479 => x"d4ff49dc",
  2480 => x"86c887e0",
  2481 => x"e8fa4873",
  2482 => x"e8fa4887",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
