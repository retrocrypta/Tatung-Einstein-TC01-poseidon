
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e0",x"ed",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"e0",x"ed",x"c2"),
    14 => (x"48",x"cc",x"db",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c6",x"e0"),
    19 => (x"72",x"1e",x"87",x"fd"),
    20 => (x"12",x"1e",x"73",x"1e"),
    21 => (x"ca",x"02",x"11",x"48"),
    22 => (x"df",x"c3",x"4b",x"87"),
    23 => (x"88",x"73",x"9b",x"98"),
    24 => (x"26",x"87",x"f0",x"02"),
    25 => (x"26",x"4a",x"26",x"4b"),
    26 => (x"1e",x"73",x"1e",x"4f"),
    27 => (x"8b",x"c1",x"1e",x"72"),
    28 => (x"12",x"87",x"ca",x"04"),
    29 => (x"c4",x"02",x"11",x"48"),
    30 => (x"f1",x"02",x"88",x"87"),
    31 => (x"26",x"4a",x"26",x"87"),
    32 => (x"1e",x"4f",x"26",x"4b"),
    33 => (x"1e",x"73",x"1e",x"74"),
    34 => (x"8b",x"c1",x"1e",x"72"),
    35 => (x"12",x"87",x"d0",x"04"),
    36 => (x"ca",x"02",x"11",x"48"),
    37 => (x"df",x"c3",x"4c",x"87"),
    38 => (x"88",x"74",x"9c",x"98"),
    39 => (x"26",x"87",x"eb",x"02"),
    40 => (x"26",x"4b",x"26",x"4a"),
    41 => (x"1e",x"4f",x"26",x"4c"),
    42 => (x"73",x"81",x"48",x"73"),
    43 => (x"87",x"c5",x"02",x"a9"),
    44 => (x"f6",x"05",x"53",x"12"),
    45 => (x"1e",x"4f",x"26",x"87"),
    46 => (x"66",x"c4",x"4a",x"71"),
    47 => (x"88",x"c1",x"48",x"49"),
    48 => (x"71",x"58",x"a6",x"c8"),
    49 => (x"87",x"d4",x"02",x"99"),
    50 => (x"d4",x"ff",x"48",x"12"),
    51 => (x"66",x"c4",x"78",x"08"),
    52 => (x"88",x"c1",x"48",x"49"),
    53 => (x"71",x"58",x"a6",x"c8"),
    54 => (x"87",x"ec",x"05",x"99"),
    55 => (x"71",x"1e",x"4f",x"26"),
    56 => (x"49",x"66",x"c4",x"4a"),
    57 => (x"c8",x"88",x"c1",x"48"),
    58 => (x"99",x"71",x"58",x"a6"),
    59 => (x"ff",x"87",x"d6",x"02"),
    60 => (x"ff",x"c3",x"48",x"d4"),
    61 => (x"c4",x"52",x"68",x"78"),
    62 => (x"c1",x"48",x"49",x"66"),
    63 => (x"58",x"a6",x"c8",x"88"),
    64 => (x"ea",x"05",x"99",x"71"),
    65 => (x"1e",x"4f",x"26",x"87"),
    66 => (x"d4",x"ff",x"1e",x"73"),
    67 => (x"7b",x"ff",x"c3",x"4b"),
    68 => (x"ff",x"c3",x"4a",x"6b"),
    69 => (x"c8",x"49",x"6b",x"7b"),
    70 => (x"c3",x"b1",x"72",x"32"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"b2",x"71",x"31",x"c8"),
    73 => (x"6b",x"7b",x"ff",x"c3"),
    74 => (x"72",x"32",x"c8",x"49"),
    75 => (x"c4",x"48",x"71",x"b1"),
    76 => (x"26",x"4d",x"26",x"87"),
    77 => (x"26",x"4b",x"26",x"4c"),
    78 => (x"5b",x"5e",x"0e",x"4f"),
    79 => (x"71",x"0e",x"5d",x"5c"),
    80 => (x"4c",x"d4",x"ff",x"4a"),
    81 => (x"ff",x"c3",x"48",x"72"),
    82 => (x"c2",x"7c",x"70",x"98"),
    83 => (x"05",x"bf",x"cc",x"db"),
    84 => (x"66",x"d0",x"87",x"c8"),
    85 => (x"d4",x"30",x"c9",x"48"),
    86 => (x"66",x"d0",x"58",x"a6"),
    87 => (x"71",x"29",x"d8",x"49"),
    88 => (x"98",x"ff",x"c3",x"48"),
    89 => (x"66",x"d0",x"7c",x"70"),
    90 => (x"71",x"29",x"d0",x"49"),
    91 => (x"98",x"ff",x"c3",x"48"),
    92 => (x"66",x"d0",x"7c",x"70"),
    93 => (x"71",x"29",x"c8",x"49"),
    94 => (x"98",x"ff",x"c3",x"48"),
    95 => (x"66",x"d0",x"7c",x"70"),
    96 => (x"98",x"ff",x"c3",x"48"),
    97 => (x"49",x"72",x"7c",x"70"),
    98 => (x"48",x"71",x"29",x"d0"),
    99 => (x"70",x"98",x"ff",x"c3"),
   100 => (x"c9",x"4b",x"6c",x"7c"),
   101 => (x"c3",x"4d",x"ff",x"f0"),
   102 => (x"d0",x"05",x"ab",x"ff"),
   103 => (x"7c",x"ff",x"c3",x"87"),
   104 => (x"8d",x"c1",x"4b",x"6c"),
   105 => (x"c3",x"87",x"c6",x"02"),
   106 => (x"f0",x"02",x"ab",x"ff"),
   107 => (x"fd",x"48",x"73",x"87"),
   108 => (x"c0",x"1e",x"87",x"ff"),
   109 => (x"48",x"d4",x"ff",x"49"),
   110 => (x"c1",x"78",x"ff",x"c3"),
   111 => (x"b7",x"c8",x"c3",x"81"),
   112 => (x"87",x"f1",x"04",x"a9"),
   113 => (x"73",x"1e",x"4f",x"26"),
   114 => (x"c4",x"87",x"e7",x"1e"),
   115 => (x"c0",x"4b",x"df",x"f8"),
   116 => (x"f0",x"ff",x"c0",x"1e"),
   117 => (x"fd",x"49",x"f7",x"c1"),
   118 => (x"86",x"c4",x"87",x"df"),
   119 => (x"c0",x"05",x"a8",x"c1"),
   120 => (x"d4",x"ff",x"87",x"ea"),
   121 => (x"78",x"ff",x"c3",x"48"),
   122 => (x"c0",x"c0",x"c0",x"c1"),
   123 => (x"c0",x"1e",x"c0",x"c0"),
   124 => (x"e9",x"c1",x"f0",x"e1"),
   125 => (x"87",x"c1",x"fd",x"49"),
   126 => (x"98",x"70",x"86",x"c4"),
   127 => (x"ff",x"87",x"ca",x"05"),
   128 => (x"ff",x"c3",x"48",x"d4"),
   129 => (x"cb",x"48",x"c1",x"78"),
   130 => (x"87",x"e6",x"fe",x"87"),
   131 => (x"fe",x"05",x"8b",x"c1"),
   132 => (x"48",x"c0",x"87",x"fd"),
   133 => (x"1e",x"87",x"de",x"fc"),
   134 => (x"d4",x"ff",x"1e",x"73"),
   135 => (x"78",x"ff",x"c3",x"48"),
   136 => (x"1e",x"c0",x"4b",x"d3"),
   137 => (x"c1",x"f0",x"ff",x"c0"),
   138 => (x"cc",x"fc",x"49",x"c1"),
   139 => (x"70",x"86",x"c4",x"87"),
   140 => (x"87",x"ca",x"05",x"98"),
   141 => (x"c3",x"48",x"d4",x"ff"),
   142 => (x"48",x"c1",x"78",x"ff"),
   143 => (x"f1",x"fd",x"87",x"cb"),
   144 => (x"05",x"8b",x"c1",x"87"),
   145 => (x"c0",x"87",x"db",x"ff"),
   146 => (x"87",x"e9",x"fb",x"48"),
   147 => (x"5c",x"5b",x"5e",x"0e"),
   148 => (x"4c",x"d4",x"ff",x"0e"),
   149 => (x"c6",x"87",x"db",x"fd"),
   150 => (x"e1",x"c0",x"1e",x"ea"),
   151 => (x"49",x"c8",x"c1",x"f0"),
   152 => (x"c4",x"87",x"d6",x"fb"),
   153 => (x"02",x"a8",x"c1",x"86"),
   154 => (x"ea",x"fe",x"87",x"c8"),
   155 => (x"c1",x"48",x"c0",x"87"),
   156 => (x"d2",x"fa",x"87",x"e2"),
   157 => (x"cf",x"49",x"70",x"87"),
   158 => (x"c6",x"99",x"ff",x"ff"),
   159 => (x"c8",x"02",x"a9",x"ea"),
   160 => (x"87",x"d3",x"fe",x"87"),
   161 => (x"cb",x"c1",x"48",x"c0"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"fc",x"4b",x"f1",x"c0"),
   164 => (x"98",x"70",x"87",x"f4"),
   165 => (x"87",x"eb",x"c0",x"02"),
   166 => (x"ff",x"c0",x"1e",x"c0"),
   167 => (x"49",x"fa",x"c1",x"f0"),
   168 => (x"c4",x"87",x"d6",x"fa"),
   169 => (x"05",x"98",x"70",x"86"),
   170 => (x"ff",x"c3",x"87",x"d9"),
   171 => (x"c3",x"49",x"6c",x"7c"),
   172 => (x"7c",x"7c",x"7c",x"ff"),
   173 => (x"99",x"c0",x"c1",x"7c"),
   174 => (x"c1",x"87",x"c4",x"02"),
   175 => (x"c0",x"87",x"d5",x"48"),
   176 => (x"c2",x"87",x"d1",x"48"),
   177 => (x"87",x"c4",x"05",x"ab"),
   178 => (x"87",x"c8",x"48",x"c0"),
   179 => (x"fe",x"05",x"8b",x"c1"),
   180 => (x"48",x"c0",x"87",x"fd"),
   181 => (x"1e",x"87",x"dc",x"f9"),
   182 => (x"db",x"c2",x"1e",x"73"),
   183 => (x"78",x"c1",x"48",x"cc"),
   184 => (x"d0",x"ff",x"4b",x"c7"),
   185 => (x"fb",x"78",x"c2",x"48"),
   186 => (x"d0",x"ff",x"87",x"c8"),
   187 => (x"c0",x"78",x"c3",x"48"),
   188 => (x"d0",x"e5",x"c0",x"1e"),
   189 => (x"f8",x"49",x"c0",x"c1"),
   190 => (x"86",x"c4",x"87",x"ff"),
   191 => (x"c1",x"05",x"a8",x"c1"),
   192 => (x"ab",x"c2",x"4b",x"87"),
   193 => (x"c0",x"87",x"c5",x"05"),
   194 => (x"87",x"f9",x"c0",x"48"),
   195 => (x"ff",x"05",x"8b",x"c1"),
   196 => (x"f7",x"fc",x"87",x"d0"),
   197 => (x"d0",x"db",x"c2",x"87"),
   198 => (x"05",x"98",x"70",x"58"),
   199 => (x"1e",x"c1",x"87",x"cd"),
   200 => (x"c1",x"f0",x"ff",x"c0"),
   201 => (x"d0",x"f8",x"49",x"d0"),
   202 => (x"ff",x"86",x"c4",x"87"),
   203 => (x"ff",x"c3",x"48",x"d4"),
   204 => (x"87",x"dd",x"c4",x"78"),
   205 => (x"58",x"d4",x"db",x"c2"),
   206 => (x"c2",x"48",x"d0",x"ff"),
   207 => (x"48",x"d4",x"ff",x"78"),
   208 => (x"c1",x"78",x"ff",x"c3"),
   209 => (x"87",x"ed",x"f7",x"48"),
   210 => (x"5c",x"5b",x"5e",x"0e"),
   211 => (x"4a",x"71",x"0e",x"5d"),
   212 => (x"ff",x"4d",x"ff",x"c3"),
   213 => (x"7c",x"75",x"4c",x"d4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"7c",x"75",x"78",x"c3"),
   216 => (x"ff",x"c0",x"1e",x"72"),
   217 => (x"49",x"d8",x"c1",x"f0"),
   218 => (x"c4",x"87",x"ce",x"f7"),
   219 => (x"02",x"98",x"70",x"86"),
   220 => (x"48",x"c1",x"87",x"c5"),
   221 => (x"75",x"87",x"ee",x"c0"),
   222 => (x"7c",x"fe",x"c3",x"7c"),
   223 => (x"d4",x"1e",x"c0",x"c8"),
   224 => (x"f2",x"f4",x"49",x"66"),
   225 => (x"75",x"86",x"c4",x"87"),
   226 => (x"75",x"7c",x"75",x"7c"),
   227 => (x"e0",x"da",x"d8",x"7c"),
   228 => (x"6c",x"7c",x"75",x"4b"),
   229 => (x"c1",x"87",x"c5",x"05"),
   230 => (x"87",x"f5",x"05",x"8b"),
   231 => (x"d0",x"ff",x"7c",x"75"),
   232 => (x"c0",x"78",x"c2",x"48"),
   233 => (x"87",x"c9",x"f6",x"48"),
   234 => (x"5c",x"5b",x"5e",x"0e"),
   235 => (x"4b",x"71",x"0e",x"5d"),
   236 => (x"ee",x"c5",x"4c",x"c0"),
   237 => (x"ff",x"4a",x"df",x"cd"),
   238 => (x"ff",x"c3",x"48",x"d4"),
   239 => (x"c3",x"48",x"68",x"78"),
   240 => (x"c0",x"05",x"a8",x"fe"),
   241 => (x"d4",x"ff",x"87",x"fe"),
   242 => (x"02",x"9b",x"73",x"4d"),
   243 => (x"66",x"d0",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c8"),
   246 => (x"d0",x"ff",x"87",x"d6"),
   247 => (x"78",x"d1",x"c4",x"48"),
   248 => (x"d0",x"7d",x"ff",x"c3"),
   249 => (x"88",x"c1",x"48",x"66"),
   250 => (x"70",x"58",x"a6",x"d4"),
   251 => (x"87",x"f0",x"05",x"98"),
   252 => (x"c3",x"48",x"d4",x"ff"),
   253 => (x"73",x"78",x"78",x"ff"),
   254 => (x"87",x"c5",x"05",x"9b"),
   255 => (x"d0",x"48",x"d0",x"ff"),
   256 => (x"4c",x"4a",x"c1",x"78"),
   257 => (x"fe",x"05",x"8a",x"c1"),
   258 => (x"48",x"74",x"87",x"ed"),
   259 => (x"1e",x"87",x"e2",x"f4"),
   260 => (x"4a",x"71",x"1e",x"73"),
   261 => (x"d4",x"ff",x"4b",x"c0"),
   262 => (x"78",x"ff",x"c3",x"48"),
   263 => (x"c4",x"48",x"d0",x"ff"),
   264 => (x"d4",x"ff",x"78",x"c3"),
   265 => (x"78",x"ff",x"c3",x"48"),
   266 => (x"ff",x"c0",x"1e",x"72"),
   267 => (x"49",x"d1",x"c1",x"f0"),
   268 => (x"c4",x"87",x"c6",x"f4"),
   269 => (x"05",x"98",x"70",x"86"),
   270 => (x"c0",x"c8",x"87",x"d2"),
   271 => (x"49",x"66",x"cc",x"1e"),
   272 => (x"c4",x"87",x"e5",x"fd"),
   273 => (x"ff",x"4b",x"70",x"86"),
   274 => (x"78",x"c2",x"48",x"d0"),
   275 => (x"e4",x"f3",x"48",x"73"),
   276 => (x"5b",x"5e",x"0e",x"87"),
   277 => (x"c0",x"0e",x"5d",x"5c"),
   278 => (x"f0",x"ff",x"c0",x"1e"),
   279 => (x"f3",x"49",x"c9",x"c1"),
   280 => (x"1e",x"d2",x"87",x"d7"),
   281 => (x"49",x"d4",x"db",x"c2"),
   282 => (x"c8",x"87",x"fd",x"fc"),
   283 => (x"c1",x"4c",x"c0",x"86"),
   284 => (x"ac",x"b7",x"d2",x"84"),
   285 => (x"c2",x"87",x"f8",x"04"),
   286 => (x"bf",x"97",x"d4",x"db"),
   287 => (x"99",x"c0",x"c3",x"49"),
   288 => (x"05",x"a9",x"c0",x"c1"),
   289 => (x"c2",x"87",x"e7",x"c0"),
   290 => (x"bf",x"97",x"db",x"db"),
   291 => (x"c2",x"31",x"d0",x"49"),
   292 => (x"bf",x"97",x"dc",x"db"),
   293 => (x"72",x"32",x"c8",x"4a"),
   294 => (x"dd",x"db",x"c2",x"b1"),
   295 => (x"b1",x"4a",x"bf",x"97"),
   296 => (x"ff",x"cf",x"4c",x"71"),
   297 => (x"c1",x"9c",x"ff",x"ff"),
   298 => (x"c1",x"34",x"ca",x"84"),
   299 => (x"db",x"c2",x"87",x"e7"),
   300 => (x"49",x"bf",x"97",x"dd"),
   301 => (x"99",x"c6",x"31",x"c1"),
   302 => (x"97",x"de",x"db",x"c2"),
   303 => (x"b7",x"c7",x"4a",x"bf"),
   304 => (x"c2",x"b1",x"72",x"2a"),
   305 => (x"bf",x"97",x"d9",x"db"),
   306 => (x"9d",x"cf",x"4d",x"4a"),
   307 => (x"97",x"da",x"db",x"c2"),
   308 => (x"9a",x"c3",x"4a",x"bf"),
   309 => (x"db",x"c2",x"32",x"ca"),
   310 => (x"4b",x"bf",x"97",x"db"),
   311 => (x"b2",x"73",x"33",x"c2"),
   312 => (x"97",x"dc",x"db",x"c2"),
   313 => (x"c0",x"c3",x"4b",x"bf"),
   314 => (x"2b",x"b7",x"c6",x"9b"),
   315 => (x"81",x"c2",x"b2",x"73"),
   316 => (x"30",x"71",x"48",x"c1"),
   317 => (x"48",x"c1",x"49",x"70"),
   318 => (x"4d",x"70",x"30",x"75"),
   319 => (x"84",x"c1",x"4c",x"72"),
   320 => (x"c0",x"c8",x"94",x"71"),
   321 => (x"cc",x"06",x"ad",x"b7"),
   322 => (x"b7",x"34",x"c1",x"87"),
   323 => (x"b7",x"c0",x"c8",x"2d"),
   324 => (x"f4",x"ff",x"01",x"ad"),
   325 => (x"f0",x"48",x"74",x"87"),
   326 => (x"5e",x"0e",x"87",x"d7"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"e3",x"c2",x"86",x"f8"),
   329 => (x"78",x"c0",x"48",x"fa"),
   330 => (x"1e",x"f2",x"db",x"c2"),
   331 => (x"de",x"fb",x"49",x"c0"),
   332 => (x"70",x"86",x"c4",x"87"),
   333 => (x"87",x"c5",x"05",x"98"),
   334 => (x"c0",x"c9",x"48",x"c0"),
   335 => (x"c1",x"4d",x"c0",x"87"),
   336 => (x"dd",x"f2",x"c0",x"7e"),
   337 => (x"dc",x"c2",x"49",x"bf"),
   338 => (x"c8",x"71",x"4a",x"e8"),
   339 => (x"87",x"d9",x"ec",x"4b"),
   340 => (x"c2",x"05",x"98",x"70"),
   341 => (x"c0",x"7e",x"c0",x"87"),
   342 => (x"49",x"bf",x"d9",x"f2"),
   343 => (x"4a",x"c4",x"dd",x"c2"),
   344 => (x"ec",x"4b",x"c8",x"71"),
   345 => (x"98",x"70",x"87",x"c3"),
   346 => (x"c0",x"87",x"c2",x"05"),
   347 => (x"c0",x"02",x"6e",x"7e"),
   348 => (x"e2",x"c2",x"87",x"fd"),
   349 => (x"c2",x"4d",x"bf",x"f8"),
   350 => (x"bf",x"9f",x"f0",x"e3"),
   351 => (x"d6",x"c5",x"48",x"7e"),
   352 => (x"c7",x"05",x"a8",x"ea"),
   353 => (x"f8",x"e2",x"c2",x"87"),
   354 => (x"87",x"ce",x"4d",x"bf"),
   355 => (x"e9",x"ca",x"48",x"6e"),
   356 => (x"c5",x"02",x"a8",x"d5"),
   357 => (x"c7",x"48",x"c0",x"87"),
   358 => (x"db",x"c2",x"87",x"e3"),
   359 => (x"49",x"75",x"1e",x"f2"),
   360 => (x"c4",x"87",x"ec",x"f9"),
   361 => (x"05",x"98",x"70",x"86"),
   362 => (x"48",x"c0",x"87",x"c5"),
   363 => (x"c0",x"87",x"ce",x"c7"),
   364 => (x"49",x"bf",x"d9",x"f2"),
   365 => (x"4a",x"c4",x"dd",x"c2"),
   366 => (x"ea",x"4b",x"c8",x"71"),
   367 => (x"98",x"70",x"87",x"eb"),
   368 => (x"c2",x"87",x"c8",x"05"),
   369 => (x"c1",x"48",x"fa",x"e3"),
   370 => (x"c0",x"87",x"da",x"78"),
   371 => (x"49",x"bf",x"dd",x"f2"),
   372 => (x"4a",x"e8",x"dc",x"c2"),
   373 => (x"ea",x"4b",x"c8",x"71"),
   374 => (x"98",x"70",x"87",x"cf"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"d8",x"c6",x"48",x"c0"),
   377 => (x"f0",x"e3",x"c2",x"87"),
   378 => (x"c1",x"49",x"bf",x"97"),
   379 => (x"c0",x"05",x"a9",x"d5"),
   380 => (x"e3",x"c2",x"87",x"cd"),
   381 => (x"49",x"bf",x"97",x"f1"),
   382 => (x"02",x"a9",x"ea",x"c2"),
   383 => (x"c0",x"87",x"c5",x"c0"),
   384 => (x"87",x"f9",x"c5",x"48"),
   385 => (x"97",x"f2",x"db",x"c2"),
   386 => (x"c3",x"48",x"7e",x"bf"),
   387 => (x"c0",x"02",x"a8",x"e9"),
   388 => (x"48",x"6e",x"87",x"ce"),
   389 => (x"02",x"a8",x"eb",x"c3"),
   390 => (x"c0",x"87",x"c5",x"c0"),
   391 => (x"87",x"dd",x"c5",x"48"),
   392 => (x"97",x"fd",x"db",x"c2"),
   393 => (x"05",x"99",x"49",x"bf"),
   394 => (x"c2",x"87",x"cc",x"c0"),
   395 => (x"bf",x"97",x"fe",x"db"),
   396 => (x"02",x"a9",x"c2",x"49"),
   397 => (x"c0",x"87",x"c5",x"c0"),
   398 => (x"87",x"c1",x"c5",x"48"),
   399 => (x"97",x"ff",x"db",x"c2"),
   400 => (x"e3",x"c2",x"48",x"bf"),
   401 => (x"4c",x"70",x"58",x"f6"),
   402 => (x"c2",x"88",x"c1",x"48"),
   403 => (x"c2",x"58",x"fa",x"e3"),
   404 => (x"bf",x"97",x"c0",x"dc"),
   405 => (x"c2",x"81",x"75",x"49"),
   406 => (x"bf",x"97",x"c1",x"dc"),
   407 => (x"72",x"32",x"c8",x"4a"),
   408 => (x"e8",x"c2",x"7e",x"a1"),
   409 => (x"78",x"6e",x"48",x"c7"),
   410 => (x"97",x"c2",x"dc",x"c2"),
   411 => (x"a6",x"c8",x"48",x"bf"),
   412 => (x"fa",x"e3",x"c2",x"58"),
   413 => (x"cf",x"c2",x"02",x"bf"),
   414 => (x"d9",x"f2",x"c0",x"87"),
   415 => (x"dd",x"c2",x"49",x"bf"),
   416 => (x"c8",x"71",x"4a",x"c4"),
   417 => (x"87",x"e1",x"e7",x"4b"),
   418 => (x"c0",x"02",x"98",x"70"),
   419 => (x"48",x"c0",x"87",x"c5"),
   420 => (x"c2",x"87",x"ea",x"c3"),
   421 => (x"4c",x"bf",x"f2",x"e3"),
   422 => (x"5c",x"db",x"e8",x"c2"),
   423 => (x"97",x"d7",x"dc",x"c2"),
   424 => (x"31",x"c8",x"49",x"bf"),
   425 => (x"97",x"d6",x"dc",x"c2"),
   426 => (x"49",x"a1",x"4a",x"bf"),
   427 => (x"97",x"d8",x"dc",x"c2"),
   428 => (x"32",x"d0",x"4a",x"bf"),
   429 => (x"c2",x"49",x"a1",x"72"),
   430 => (x"bf",x"97",x"d9",x"dc"),
   431 => (x"72",x"32",x"d8",x"4a"),
   432 => (x"66",x"c4",x"49",x"a1"),
   433 => (x"c7",x"e8",x"c2",x"91"),
   434 => (x"e8",x"c2",x"81",x"bf"),
   435 => (x"dc",x"c2",x"59",x"cf"),
   436 => (x"4a",x"bf",x"97",x"df"),
   437 => (x"dc",x"c2",x"32",x"c8"),
   438 => (x"4b",x"bf",x"97",x"de"),
   439 => (x"dc",x"c2",x"4a",x"a2"),
   440 => (x"4b",x"bf",x"97",x"e0"),
   441 => (x"a2",x"73",x"33",x"d0"),
   442 => (x"e1",x"dc",x"c2",x"4a"),
   443 => (x"cf",x"4b",x"bf",x"97"),
   444 => (x"73",x"33",x"d8",x"9b"),
   445 => (x"e8",x"c2",x"4a",x"a2"),
   446 => (x"8a",x"c2",x"5a",x"d3"),
   447 => (x"e8",x"c2",x"92",x"74"),
   448 => (x"a1",x"72",x"48",x"d3"),
   449 => (x"87",x"c1",x"c1",x"78"),
   450 => (x"97",x"c4",x"dc",x"c2"),
   451 => (x"31",x"c8",x"49",x"bf"),
   452 => (x"97",x"c3",x"dc",x"c2"),
   453 => (x"49",x"a1",x"4a",x"bf"),
   454 => (x"ff",x"c7",x"31",x"c5"),
   455 => (x"c2",x"29",x"c9",x"81"),
   456 => (x"c2",x"59",x"db",x"e8"),
   457 => (x"bf",x"97",x"c9",x"dc"),
   458 => (x"c2",x"32",x"c8",x"4a"),
   459 => (x"bf",x"97",x"c8",x"dc"),
   460 => (x"c4",x"4a",x"a2",x"4b"),
   461 => (x"82",x"6e",x"92",x"66"),
   462 => (x"5a",x"d7",x"e8",x"c2"),
   463 => (x"48",x"cf",x"e8",x"c2"),
   464 => (x"e8",x"c2",x"78",x"c0"),
   465 => (x"a1",x"72",x"48",x"cb"),
   466 => (x"db",x"e8",x"c2",x"78"),
   467 => (x"cf",x"e8",x"c2",x"48"),
   468 => (x"e8",x"c2",x"78",x"bf"),
   469 => (x"e8",x"c2",x"48",x"df"),
   470 => (x"c2",x"78",x"bf",x"d3"),
   471 => (x"02",x"bf",x"fa",x"e3"),
   472 => (x"74",x"87",x"c9",x"c0"),
   473 => (x"70",x"30",x"c4",x"48"),
   474 => (x"87",x"c9",x"c0",x"7e"),
   475 => (x"bf",x"d7",x"e8",x"c2"),
   476 => (x"70",x"30",x"c4",x"48"),
   477 => (x"fe",x"e3",x"c2",x"7e"),
   478 => (x"c1",x"78",x"6e",x"48"),
   479 => (x"26",x"8e",x"f8",x"48"),
   480 => (x"26",x"4c",x"26",x"4d"),
   481 => (x"0e",x"4f",x"26",x"4b"),
   482 => (x"5d",x"5c",x"5b",x"5e"),
   483 => (x"c2",x"4a",x"71",x"0e"),
   484 => (x"02",x"bf",x"fa",x"e3"),
   485 => (x"4b",x"72",x"87",x"cb"),
   486 => (x"4d",x"72",x"2b",x"c7"),
   487 => (x"c9",x"9d",x"ff",x"c1"),
   488 => (x"c8",x"4b",x"72",x"87"),
   489 => (x"c3",x"4d",x"72",x"2b"),
   490 => (x"e8",x"c2",x"9d",x"ff"),
   491 => (x"c0",x"83",x"bf",x"c7"),
   492 => (x"ab",x"bf",x"d5",x"f2"),
   493 => (x"c0",x"87",x"d9",x"02"),
   494 => (x"c2",x"5b",x"d9",x"f2"),
   495 => (x"73",x"1e",x"f2",x"db"),
   496 => (x"87",x"cb",x"f1",x"49"),
   497 => (x"98",x"70",x"86",x"c4"),
   498 => (x"c0",x"87",x"c5",x"05"),
   499 => (x"87",x"e6",x"c0",x"48"),
   500 => (x"bf",x"fa",x"e3",x"c2"),
   501 => (x"75",x"87",x"d2",x"02"),
   502 => (x"c2",x"91",x"c4",x"49"),
   503 => (x"69",x"81",x"f2",x"db"),
   504 => (x"ff",x"ff",x"cf",x"4c"),
   505 => (x"cb",x"9c",x"ff",x"ff"),
   506 => (x"c2",x"49",x"75",x"87"),
   507 => (x"f2",x"db",x"c2",x"91"),
   508 => (x"4c",x"69",x"9f",x"81"),
   509 => (x"c6",x"fe",x"48",x"74"),
   510 => (x"5b",x"5e",x"0e",x"87"),
   511 => (x"f8",x"0e",x"5d",x"5c"),
   512 => (x"9c",x"4c",x"71",x"86"),
   513 => (x"c0",x"87",x"c5",x"05"),
   514 => (x"87",x"c0",x"c3",x"48"),
   515 => (x"48",x"7e",x"a4",x"c8"),
   516 => (x"66",x"d8",x"78",x"c0"),
   517 => (x"d8",x"87",x"c7",x"02"),
   518 => (x"05",x"bf",x"97",x"66"),
   519 => (x"48",x"c0",x"87",x"c5"),
   520 => (x"c0",x"87",x"e9",x"c2"),
   521 => (x"49",x"49",x"c1",x"1e"),
   522 => (x"c4",x"87",x"d3",x"ca"),
   523 => (x"9d",x"4d",x"70",x"86"),
   524 => (x"87",x"c2",x"c1",x"02"),
   525 => (x"4a",x"c2",x"e4",x"c2"),
   526 => (x"e0",x"49",x"66",x"d8"),
   527 => (x"98",x"70",x"87",x"d0"),
   528 => (x"87",x"f2",x"c0",x"02"),
   529 => (x"66",x"d8",x"4a",x"75"),
   530 => (x"e0",x"4b",x"cb",x"49"),
   531 => (x"98",x"70",x"87",x"f5"),
   532 => (x"87",x"e2",x"c0",x"02"),
   533 => (x"9d",x"75",x"1e",x"c0"),
   534 => (x"c8",x"87",x"c7",x"02"),
   535 => (x"78",x"c0",x"48",x"a6"),
   536 => (x"a6",x"c8",x"87",x"c5"),
   537 => (x"c8",x"78",x"c1",x"48"),
   538 => (x"d1",x"c9",x"49",x"66"),
   539 => (x"70",x"86",x"c4",x"87"),
   540 => (x"fe",x"05",x"9d",x"4d"),
   541 => (x"9d",x"75",x"87",x"fe"),
   542 => (x"87",x"ce",x"c1",x"02"),
   543 => (x"6e",x"49",x"a5",x"dc"),
   544 => (x"da",x"78",x"69",x"48"),
   545 => (x"a6",x"c4",x"49",x"a5"),
   546 => (x"78",x"a4",x"c4",x"48"),
   547 => (x"c4",x"48",x"69",x"9f"),
   548 => (x"c2",x"78",x"08",x"66"),
   549 => (x"02",x"bf",x"fa",x"e3"),
   550 => (x"a5",x"d4",x"87",x"d2"),
   551 => (x"49",x"69",x"9f",x"49"),
   552 => (x"99",x"ff",x"ff",x"c0"),
   553 => (x"30",x"d0",x"48",x"71"),
   554 => (x"87",x"c2",x"7e",x"70"),
   555 => (x"48",x"6e",x"7e",x"c0"),
   556 => (x"80",x"bf",x"66",x"c4"),
   557 => (x"78",x"08",x"66",x"c4"),
   558 => (x"a4",x"cc",x"7c",x"c0"),
   559 => (x"bf",x"66",x"c4",x"49"),
   560 => (x"49",x"a4",x"d0",x"79"),
   561 => (x"48",x"c1",x"79",x"c0"),
   562 => (x"48",x"c0",x"87",x"c2"),
   563 => (x"ee",x"fa",x"8e",x"f8"),
   564 => (x"5b",x"5e",x"0e",x"87"),
   565 => (x"4c",x"71",x"0e",x"5c"),
   566 => (x"cb",x"c1",x"02",x"9c"),
   567 => (x"49",x"a4",x"c8",x"87"),
   568 => (x"c3",x"c1",x"02",x"69"),
   569 => (x"cc",x"49",x"6c",x"87"),
   570 => (x"80",x"71",x"48",x"66"),
   571 => (x"70",x"58",x"a6",x"d0"),
   572 => (x"f6",x"e3",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e5",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"ff",x"f9",x"49"),
   578 => (x"e3",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"f2"),
   580 => (x"cc",x"7c",x"71",x"81"),
   581 => (x"e3",x"c2",x"b9",x"66"),
   582 => (x"ff",x"4a",x"bf",x"f6"),
   583 => (x"71",x"99",x"72",x"ba"),
   584 => (x"db",x"ff",x"05",x"99"),
   585 => (x"7c",x"66",x"cc",x"87"),
   586 => (x"1e",x"87",x"d6",x"f9"),
   587 => (x"4b",x"71",x"1e",x"73"),
   588 => (x"87",x"c7",x"02",x"9b"),
   589 => (x"69",x"49",x"a3",x"c8"),
   590 => (x"c0",x"87",x"c5",x"05"),
   591 => (x"87",x"f6",x"c0",x"48"),
   592 => (x"bf",x"cb",x"e8",x"c2"),
   593 => (x"4a",x"a3",x"c4",x"49"),
   594 => (x"8a",x"c2",x"4a",x"6a"),
   595 => (x"bf",x"f2",x"e3",x"c2"),
   596 => (x"49",x"a1",x"72",x"92"),
   597 => (x"bf",x"f6",x"e3",x"c2"),
   598 => (x"72",x"9a",x"6b",x"4a"),
   599 => (x"f2",x"c0",x"49",x"a1"),
   600 => (x"66",x"c8",x"59",x"d9"),
   601 => (x"e6",x"ea",x"71",x"1e"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"87",x"c4",x"05",x"98"),
   604 => (x"87",x"c2",x"48",x"c0"),
   605 => (x"ca",x"f8",x"48",x"c1"),
   606 => (x"1e",x"73",x"1e",x"87"),
   607 => (x"02",x"9b",x"4b",x"71"),
   608 => (x"a3",x"c8",x"87",x"c7"),
   609 => (x"c5",x"05",x"69",x"49"),
   610 => (x"c0",x"48",x"c0",x"87"),
   611 => (x"e8",x"c2",x"87",x"f6"),
   612 => (x"c4",x"49",x"bf",x"cb"),
   613 => (x"4a",x"6a",x"4a",x"a3"),
   614 => (x"e3",x"c2",x"8a",x"c2"),
   615 => (x"72",x"92",x"bf",x"f2"),
   616 => (x"e3",x"c2",x"49",x"a1"),
   617 => (x"6b",x"4a",x"bf",x"f6"),
   618 => (x"49",x"a1",x"72",x"9a"),
   619 => (x"59",x"d9",x"f2",x"c0"),
   620 => (x"71",x"1e",x"66",x"c8"),
   621 => (x"c4",x"87",x"d1",x"e6"),
   622 => (x"05",x"98",x"70",x"86"),
   623 => (x"48",x"c0",x"87",x"c4"),
   624 => (x"48",x"c1",x"87",x"c2"),
   625 => (x"0e",x"87",x"fc",x"f6"),
   626 => (x"5d",x"5c",x"5b",x"5e"),
   627 => (x"4b",x"71",x"1e",x"0e"),
   628 => (x"73",x"4d",x"66",x"d4"),
   629 => (x"cc",x"c1",x"02",x"9b"),
   630 => (x"49",x"a3",x"c8",x"87"),
   631 => (x"c4",x"c1",x"02",x"69"),
   632 => (x"4c",x"a3",x"d0",x"87"),
   633 => (x"bf",x"f6",x"e3",x"c2"),
   634 => (x"6c",x"b9",x"ff",x"49"),
   635 => (x"d4",x"7e",x"99",x"4a"),
   636 => (x"cd",x"06",x"a9",x"66"),
   637 => (x"7c",x"7b",x"c0",x"87"),
   638 => (x"c4",x"4a",x"a3",x"cc"),
   639 => (x"79",x"6a",x"49",x"a3"),
   640 => (x"49",x"72",x"87",x"ca"),
   641 => (x"d4",x"99",x"c0",x"f8"),
   642 => (x"8d",x"71",x"4d",x"66"),
   643 => (x"29",x"c9",x"49",x"75"),
   644 => (x"49",x"73",x"1e",x"71"),
   645 => (x"c2",x"87",x"fa",x"fa"),
   646 => (x"73",x"1e",x"f2",x"db"),
   647 => (x"87",x"cb",x"fc",x"49"),
   648 => (x"66",x"d4",x"86",x"c8"),
   649 => (x"d6",x"f5",x"26",x"7c"),
   650 => (x"1e",x"73",x"1e",x"87"),
   651 => (x"02",x"9b",x"4b",x"71"),
   652 => (x"c2",x"87",x"e4",x"c0"),
   653 => (x"73",x"5b",x"df",x"e8"),
   654 => (x"c2",x"8a",x"c2",x"4a"),
   655 => (x"49",x"bf",x"f2",x"e3"),
   656 => (x"cb",x"e8",x"c2",x"92"),
   657 => (x"80",x"72",x"48",x"bf"),
   658 => (x"58",x"e3",x"e8",x"c2"),
   659 => (x"30",x"c4",x"48",x"71"),
   660 => (x"58",x"c2",x"e4",x"c2"),
   661 => (x"c2",x"87",x"ed",x"c0"),
   662 => (x"c2",x"48",x"db",x"e8"),
   663 => (x"78",x"bf",x"cf",x"e8"),
   664 => (x"48",x"df",x"e8",x"c2"),
   665 => (x"bf",x"d3",x"e8",x"c2"),
   666 => (x"fa",x"e3",x"c2",x"78"),
   667 => (x"87",x"c9",x"02",x"bf"),
   668 => (x"bf",x"f2",x"e3",x"c2"),
   669 => (x"c7",x"31",x"c4",x"49"),
   670 => (x"d7",x"e8",x"c2",x"87"),
   671 => (x"31",x"c4",x"49",x"bf"),
   672 => (x"59",x"c2",x"e4",x"c2"),
   673 => (x"0e",x"87",x"fc",x"f3"),
   674 => (x"0e",x"5c",x"5b",x"5e"),
   675 => (x"4b",x"c0",x"4a",x"71"),
   676 => (x"c0",x"02",x"9a",x"72"),
   677 => (x"a2",x"da",x"87",x"e0"),
   678 => (x"4b",x"69",x"9f",x"49"),
   679 => (x"bf",x"fa",x"e3",x"c2"),
   680 => (x"d4",x"87",x"cf",x"02"),
   681 => (x"69",x"9f",x"49",x"a2"),
   682 => (x"ff",x"c0",x"4c",x"49"),
   683 => (x"34",x"d0",x"9c",x"ff"),
   684 => (x"4c",x"c0",x"87",x"c2"),
   685 => (x"49",x"73",x"b3",x"74"),
   686 => (x"f3",x"87",x"ee",x"fd"),
   687 => (x"5e",x"0e",x"87",x"c3"),
   688 => (x"0e",x"5d",x"5c",x"5b"),
   689 => (x"4a",x"71",x"86",x"f4"),
   690 => (x"9a",x"72",x"7e",x"c0"),
   691 => (x"c2",x"87",x"d8",x"02"),
   692 => (x"c0",x"48",x"ee",x"db"),
   693 => (x"e6",x"db",x"c2",x"78"),
   694 => (x"df",x"e8",x"c2",x"48"),
   695 => (x"db",x"c2",x"78",x"bf"),
   696 => (x"e8",x"c2",x"48",x"ea"),
   697 => (x"c2",x"78",x"bf",x"db"),
   698 => (x"c0",x"48",x"cf",x"e4"),
   699 => (x"fe",x"e3",x"c2",x"50"),
   700 => (x"db",x"c2",x"49",x"bf"),
   701 => (x"71",x"4a",x"bf",x"ee"),
   702 => (x"c9",x"c4",x"03",x"aa"),
   703 => (x"cf",x"49",x"72",x"87"),
   704 => (x"e9",x"c0",x"05",x"99"),
   705 => (x"d5",x"f2",x"c0",x"87"),
   706 => (x"e6",x"db",x"c2",x"48"),
   707 => (x"db",x"c2",x"78",x"bf"),
   708 => (x"db",x"c2",x"1e",x"f2"),
   709 => (x"c2",x"49",x"bf",x"e6"),
   710 => (x"c1",x"48",x"e6",x"db"),
   711 => (x"e3",x"71",x"78",x"a1"),
   712 => (x"86",x"c4",x"87",x"ed"),
   713 => (x"48",x"d1",x"f2",x"c0"),
   714 => (x"78",x"f2",x"db",x"c2"),
   715 => (x"f2",x"c0",x"87",x"cc"),
   716 => (x"c0",x"48",x"bf",x"d1"),
   717 => (x"f2",x"c0",x"80",x"e0"),
   718 => (x"db",x"c2",x"58",x"d5"),
   719 => (x"c1",x"48",x"bf",x"ee"),
   720 => (x"f2",x"db",x"c2",x"80"),
   721 => (x"0c",x"91",x"27",x"58"),
   722 => (x"97",x"bf",x"00",x"00"),
   723 => (x"02",x"9d",x"4d",x"bf"),
   724 => (x"c3",x"87",x"e3",x"c2"),
   725 => (x"c2",x"02",x"ad",x"e5"),
   726 => (x"f2",x"c0",x"87",x"dc"),
   727 => (x"cb",x"4b",x"bf",x"d1"),
   728 => (x"4c",x"11",x"49",x"a3"),
   729 => (x"c1",x"05",x"ac",x"cf"),
   730 => (x"49",x"75",x"87",x"d2"),
   731 => (x"89",x"c1",x"99",x"df"),
   732 => (x"e4",x"c2",x"91",x"cd"),
   733 => (x"a3",x"c1",x"81",x"c2"),
   734 => (x"c3",x"51",x"12",x"4a"),
   735 => (x"51",x"12",x"4a",x"a3"),
   736 => (x"12",x"4a",x"a3",x"c5"),
   737 => (x"4a",x"a3",x"c7",x"51"),
   738 => (x"a3",x"c9",x"51",x"12"),
   739 => (x"ce",x"51",x"12",x"4a"),
   740 => (x"51",x"12",x"4a",x"a3"),
   741 => (x"12",x"4a",x"a3",x"d0"),
   742 => (x"4a",x"a3",x"d2",x"51"),
   743 => (x"a3",x"d4",x"51",x"12"),
   744 => (x"d6",x"51",x"12",x"4a"),
   745 => (x"51",x"12",x"4a",x"a3"),
   746 => (x"12",x"4a",x"a3",x"d8"),
   747 => (x"4a",x"a3",x"dc",x"51"),
   748 => (x"a3",x"de",x"51",x"12"),
   749 => (x"c1",x"51",x"12",x"4a"),
   750 => (x"87",x"fa",x"c0",x"7e"),
   751 => (x"99",x"c8",x"49",x"74"),
   752 => (x"87",x"eb",x"c0",x"05"),
   753 => (x"99",x"d0",x"49",x"74"),
   754 => (x"dc",x"87",x"d1",x"05"),
   755 => (x"cb",x"c0",x"02",x"66"),
   756 => (x"dc",x"49",x"73",x"87"),
   757 => (x"98",x"70",x"0f",x"66"),
   758 => (x"87",x"d3",x"c0",x"02"),
   759 => (x"c6",x"c0",x"05",x"6e"),
   760 => (x"c2",x"e4",x"c2",x"87"),
   761 => (x"c0",x"50",x"c0",x"48"),
   762 => (x"48",x"bf",x"d1",x"f2"),
   763 => (x"c2",x"87",x"dd",x"c2"),
   764 => (x"c0",x"48",x"cf",x"e4"),
   765 => (x"e3",x"c2",x"7e",x"50"),
   766 => (x"c2",x"49",x"bf",x"fe"),
   767 => (x"4a",x"bf",x"ee",x"db"),
   768 => (x"fb",x"04",x"aa",x"71"),
   769 => (x"e8",x"c2",x"87",x"f7"),
   770 => (x"c0",x"05",x"bf",x"df"),
   771 => (x"e3",x"c2",x"87",x"c8"),
   772 => (x"c1",x"02",x"bf",x"fa"),
   773 => (x"db",x"c2",x"87",x"f4"),
   774 => (x"ed",x"49",x"bf",x"ea"),
   775 => (x"db",x"c2",x"87",x"e9"),
   776 => (x"a6",x"c4",x"58",x"ee"),
   777 => (x"ea",x"db",x"c2",x"48"),
   778 => (x"e3",x"c2",x"78",x"bf"),
   779 => (x"c0",x"02",x"bf",x"fa"),
   780 => (x"66",x"c4",x"87",x"d8"),
   781 => (x"ff",x"ff",x"cf",x"49"),
   782 => (x"a9",x"99",x"f8",x"ff"),
   783 => (x"87",x"c5",x"c0",x"02"),
   784 => (x"e1",x"c0",x"4c",x"c0"),
   785 => (x"c0",x"4c",x"c1",x"87"),
   786 => (x"66",x"c4",x"87",x"dc"),
   787 => (x"f8",x"ff",x"cf",x"49"),
   788 => (x"c0",x"02",x"a9",x"99"),
   789 => (x"a6",x"c8",x"87",x"c8"),
   790 => (x"c0",x"78",x"c0",x"48"),
   791 => (x"a6",x"c8",x"87",x"c5"),
   792 => (x"c8",x"78",x"c1",x"48"),
   793 => (x"9c",x"74",x"4c",x"66"),
   794 => (x"87",x"de",x"c0",x"05"),
   795 => (x"c2",x"49",x"66",x"c4"),
   796 => (x"f2",x"e3",x"c2",x"89"),
   797 => (x"e8",x"c2",x"91",x"bf"),
   798 => (x"71",x"48",x"bf",x"cb"),
   799 => (x"ea",x"db",x"c2",x"80"),
   800 => (x"ee",x"db",x"c2",x"58"),
   801 => (x"f9",x"78",x"c0",x"48"),
   802 => (x"48",x"c0",x"87",x"e3"),
   803 => (x"ee",x"eb",x"8e",x"f4"),
   804 => (x"00",x"00",x"00",x"87"),
   805 => (x"ff",x"ff",x"ff",x"00"),
   806 => (x"00",x"0c",x"a1",x"ff"),
   807 => (x"00",x"0c",x"aa",x"00"),
   808 => (x"54",x"41",x"46",x"00"),
   809 => (x"20",x"20",x"32",x"33"),
   810 => (x"41",x"46",x"00",x"20"),
   811 => (x"20",x"36",x"31",x"54"),
   812 => (x"1e",x"00",x"20",x"20"),
   813 => (x"c3",x"48",x"d4",x"ff"),
   814 => (x"48",x"68",x"78",x"ff"),
   815 => (x"ff",x"1e",x"4f",x"26"),
   816 => (x"ff",x"c3",x"48",x"d4"),
   817 => (x"48",x"d0",x"ff",x"78"),
   818 => (x"ff",x"78",x"e1",x"c0"),
   819 => (x"78",x"d4",x"48",x"d4"),
   820 => (x"48",x"e3",x"e8",x"c2"),
   821 => (x"50",x"bf",x"d4",x"ff"),
   822 => (x"ff",x"1e",x"4f",x"26"),
   823 => (x"e0",x"c0",x"48",x"d0"),
   824 => (x"1e",x"4f",x"26",x"78"),
   825 => (x"70",x"87",x"cc",x"ff"),
   826 => (x"c6",x"02",x"99",x"49"),
   827 => (x"a9",x"fb",x"c0",x"87"),
   828 => (x"71",x"87",x"f1",x"05"),
   829 => (x"0e",x"4f",x"26",x"48"),
   830 => (x"0e",x"5c",x"5b",x"5e"),
   831 => (x"4c",x"c0",x"4b",x"71"),
   832 => (x"70",x"87",x"f0",x"fe"),
   833 => (x"c0",x"02",x"99",x"49"),
   834 => (x"ec",x"c0",x"87",x"f9"),
   835 => (x"f2",x"c0",x"02",x"a9"),
   836 => (x"a9",x"fb",x"c0",x"87"),
   837 => (x"87",x"eb",x"c0",x"02"),
   838 => (x"ac",x"b7",x"66",x"cc"),
   839 => (x"d0",x"87",x"c7",x"03"),
   840 => (x"87",x"c2",x"02",x"66"),
   841 => (x"99",x"71",x"53",x"71"),
   842 => (x"c1",x"87",x"c2",x"02"),
   843 => (x"87",x"c3",x"fe",x"84"),
   844 => (x"02",x"99",x"49",x"70"),
   845 => (x"ec",x"c0",x"87",x"cd"),
   846 => (x"87",x"c7",x"02",x"a9"),
   847 => (x"05",x"a9",x"fb",x"c0"),
   848 => (x"d0",x"87",x"d5",x"ff"),
   849 => (x"87",x"c3",x"02",x"66"),
   850 => (x"c0",x"7b",x"97",x"c0"),
   851 => (x"c4",x"05",x"a9",x"ec"),
   852 => (x"c5",x"4a",x"74",x"87"),
   853 => (x"c0",x"4a",x"74",x"87"),
   854 => (x"48",x"72",x"8a",x"0a"),
   855 => (x"4d",x"26",x"87",x"c2"),
   856 => (x"4b",x"26",x"4c",x"26"),
   857 => (x"fd",x"1e",x"4f",x"26"),
   858 => (x"49",x"70",x"87",x"c9"),
   859 => (x"aa",x"f0",x"c0",x"4a"),
   860 => (x"c0",x"87",x"c9",x"04"),
   861 => (x"c3",x"01",x"aa",x"f9"),
   862 => (x"8a",x"f0",x"c0",x"87"),
   863 => (x"04",x"aa",x"c1",x"c1"),
   864 => (x"da",x"c1",x"87",x"c9"),
   865 => (x"87",x"c3",x"01",x"aa"),
   866 => (x"72",x"8a",x"f7",x"c0"),
   867 => (x"0e",x"4f",x"26",x"48"),
   868 => (x"5d",x"5c",x"5b",x"5e"),
   869 => (x"71",x"86",x"f8",x"0e"),
   870 => (x"fc",x"4d",x"c0",x"4c"),
   871 => (x"4b",x"c0",x"87",x"e0"),
   872 => (x"97",x"ee",x"f8",x"c0"),
   873 => (x"a9",x"c0",x"49",x"bf"),
   874 => (x"fc",x"87",x"cf",x"04"),
   875 => (x"83",x"c1",x"87",x"f5"),
   876 => (x"97",x"ee",x"f8",x"c0"),
   877 => (x"06",x"ab",x"49",x"bf"),
   878 => (x"f8",x"c0",x"87",x"f1"),
   879 => (x"02",x"bf",x"97",x"ee"),
   880 => (x"ee",x"fb",x"87",x"cf"),
   881 => (x"99",x"49",x"70",x"87"),
   882 => (x"c0",x"87",x"c6",x"02"),
   883 => (x"f1",x"05",x"a9",x"ec"),
   884 => (x"fb",x"4b",x"c0",x"87"),
   885 => (x"7e",x"70",x"87",x"dd"),
   886 => (x"c8",x"87",x"d8",x"fb"),
   887 => (x"d2",x"fb",x"58",x"a6"),
   888 => (x"c1",x"4a",x"70",x"87"),
   889 => (x"49",x"a4",x"c8",x"83"),
   890 => (x"6e",x"49",x"69",x"97"),
   891 => (x"87",x"da",x"05",x"a9"),
   892 => (x"97",x"49",x"a4",x"c9"),
   893 => (x"66",x"c4",x"49",x"69"),
   894 => (x"87",x"ce",x"05",x"a9"),
   895 => (x"97",x"49",x"a4",x"ca"),
   896 => (x"05",x"aa",x"49",x"69"),
   897 => (x"4d",x"c1",x"87",x"c4"),
   898 => (x"48",x"6e",x"87",x"d4"),
   899 => (x"02",x"a8",x"ec",x"c0"),
   900 => (x"48",x"6e",x"87",x"c8"),
   901 => (x"05",x"a8",x"fb",x"c0"),
   902 => (x"4b",x"c0",x"87",x"c4"),
   903 => (x"9d",x"75",x"4d",x"c1"),
   904 => (x"87",x"ef",x"fe",x"02"),
   905 => (x"73",x"87",x"f3",x"fa"),
   906 => (x"fc",x"8e",x"f8",x"48"),
   907 => (x"0e",x"00",x"87",x"f0"),
   908 => (x"5d",x"5c",x"5b",x"5e"),
   909 => (x"71",x"86",x"f8",x"0e"),
   910 => (x"4b",x"d4",x"ff",x"7e"),
   911 => (x"e8",x"c2",x"1e",x"6e"),
   912 => (x"f4",x"e6",x"49",x"e8"),
   913 => (x"70",x"86",x"c4",x"87"),
   914 => (x"ea",x"c4",x"02",x"98"),
   915 => (x"d5",x"e3",x"c1",x"87"),
   916 => (x"49",x"6e",x"4d",x"bf"),
   917 => (x"c8",x"87",x"f8",x"fc"),
   918 => (x"98",x"70",x"58",x"a6"),
   919 => (x"c4",x"87",x"c5",x"05"),
   920 => (x"78",x"c1",x"48",x"a6"),
   921 => (x"c5",x"48",x"d0",x"ff"),
   922 => (x"7b",x"d5",x"c1",x"78"),
   923 => (x"c1",x"49",x"66",x"c4"),
   924 => (x"c1",x"31",x"c6",x"89"),
   925 => (x"bf",x"97",x"d3",x"e3"),
   926 => (x"b0",x"71",x"48",x"4a"),
   927 => (x"d0",x"ff",x"7b",x"70"),
   928 => (x"c2",x"78",x"c4",x"48"),
   929 => (x"bf",x"97",x"e3",x"e8"),
   930 => (x"02",x"99",x"d0",x"49"),
   931 => (x"78",x"c5",x"87",x"d7"),
   932 => (x"c0",x"7b",x"d6",x"c1"),
   933 => (x"7b",x"ff",x"c3",x"4a"),
   934 => (x"e0",x"c0",x"82",x"c1"),
   935 => (x"87",x"f5",x"04",x"aa"),
   936 => (x"c4",x"48",x"d0",x"ff"),
   937 => (x"7b",x"ff",x"c3",x"78"),
   938 => (x"c5",x"48",x"d0",x"ff"),
   939 => (x"7b",x"d3",x"c1",x"78"),
   940 => (x"78",x"c4",x"7b",x"c1"),
   941 => (x"06",x"ad",x"b7",x"c0"),
   942 => (x"c2",x"87",x"eb",x"c2"),
   943 => (x"4c",x"bf",x"f0",x"e8"),
   944 => (x"c2",x"02",x"9c",x"8d"),
   945 => (x"db",x"c2",x"87",x"c2"),
   946 => (x"a6",x"c4",x"7e",x"f2"),
   947 => (x"78",x"c0",x"c8",x"48"),
   948 => (x"ac",x"b7",x"c0",x"8c"),
   949 => (x"c8",x"87",x"c6",x"03"),
   950 => (x"c0",x"78",x"a4",x"c0"),
   951 => (x"e3",x"e8",x"c2",x"4c"),
   952 => (x"d0",x"49",x"bf",x"97"),
   953 => (x"87",x"d0",x"02",x"99"),
   954 => (x"e8",x"c2",x"1e",x"c0"),
   955 => (x"fa",x"e8",x"49",x"e8"),
   956 => (x"70",x"86",x"c4",x"87"),
   957 => (x"87",x"f5",x"c0",x"4a"),
   958 => (x"1e",x"f2",x"db",x"c2"),
   959 => (x"49",x"e8",x"e8",x"c2"),
   960 => (x"c4",x"87",x"e8",x"e8"),
   961 => (x"ff",x"4a",x"70",x"86"),
   962 => (x"c5",x"c8",x"48",x"d0"),
   963 => (x"7b",x"d4",x"c1",x"78"),
   964 => (x"7b",x"bf",x"97",x"6e"),
   965 => (x"80",x"c1",x"48",x"6e"),
   966 => (x"66",x"c4",x"7e",x"70"),
   967 => (x"c8",x"88",x"c1",x"48"),
   968 => (x"98",x"70",x"58",x"a6"),
   969 => (x"87",x"e8",x"ff",x"05"),
   970 => (x"c4",x"48",x"d0",x"ff"),
   971 => (x"05",x"9a",x"72",x"78"),
   972 => (x"48",x"c0",x"87",x"c5"),
   973 => (x"c1",x"87",x"c2",x"c1"),
   974 => (x"e8",x"e8",x"c2",x"1e"),
   975 => (x"87",x"d1",x"e6",x"49"),
   976 => (x"9c",x"74",x"86",x"c4"),
   977 => (x"87",x"fe",x"fd",x"05"),
   978 => (x"06",x"ad",x"b7",x"c0"),
   979 => (x"e8",x"c2",x"87",x"d1"),
   980 => (x"78",x"c0",x"48",x"e8"),
   981 => (x"78",x"c0",x"80",x"d0"),
   982 => (x"e8",x"c2",x"80",x"f4"),
   983 => (x"c0",x"78",x"bf",x"f4"),
   984 => (x"fd",x"01",x"ad",x"b7"),
   985 => (x"d0",x"ff",x"87",x"d5"),
   986 => (x"c1",x"78",x"c5",x"48"),
   987 => (x"7b",x"c0",x"7b",x"d3"),
   988 => (x"48",x"c1",x"78",x"c4"),
   989 => (x"c0",x"87",x"c2",x"c0"),
   990 => (x"26",x"8e",x"f8",x"48"),
   991 => (x"26",x"4c",x"26",x"4d"),
   992 => (x"0e",x"4f",x"26",x"4b"),
   993 => (x"5d",x"5c",x"5b",x"5e"),
   994 => (x"4b",x"71",x"1e",x"0e"),
   995 => (x"ab",x"4d",x"4c",x"c0"),
   996 => (x"87",x"e8",x"c0",x"04"),
   997 => (x"1e",x"cf",x"f6",x"c0"),
   998 => (x"c4",x"02",x"9d",x"75"),
   999 => (x"c2",x"4a",x"c0",x"87"),
  1000 => (x"72",x"4a",x"c1",x"87"),
  1001 => (x"87",x"d6",x"ec",x"49"),
  1002 => (x"7e",x"70",x"86",x"c4"),
  1003 => (x"05",x"6e",x"84",x"c1"),
  1004 => (x"4c",x"73",x"87",x"c2"),
  1005 => (x"ac",x"73",x"85",x"c1"),
  1006 => (x"87",x"d8",x"ff",x"06"),
  1007 => (x"fe",x"26",x"48",x"6e"),
  1008 => (x"5e",x"0e",x"87",x"f9"),
  1009 => (x"71",x"0e",x"5c",x"5b"),
  1010 => (x"02",x"66",x"cc",x"4b"),
  1011 => (x"c0",x"4c",x"87",x"d8"),
  1012 => (x"d8",x"02",x"8c",x"f0"),
  1013 => (x"c1",x"4a",x"74",x"87"),
  1014 => (x"87",x"d1",x"02",x"8a"),
  1015 => (x"87",x"cd",x"02",x"8a"),
  1016 => (x"87",x"c9",x"02",x"8a"),
  1017 => (x"49",x"73",x"87",x"d9"),
  1018 => (x"d2",x"87",x"c4",x"f9"),
  1019 => (x"c0",x"1e",x"74",x"87"),
  1020 => (x"d7",x"d9",x"c1",x"49"),
  1021 => (x"73",x"1e",x"74",x"87"),
  1022 => (x"cf",x"d9",x"c1",x"49"),
  1023 => (x"fd",x"86",x"c8",x"87"),
  1024 => (x"5e",x"0e",x"87",x"fb"),
  1025 => (x"0e",x"5d",x"5c",x"5b"),
  1026 => (x"49",x"4c",x"71",x"1e"),
  1027 => (x"e9",x"c2",x"91",x"de"),
  1028 => (x"85",x"71",x"4d",x"d0"),
  1029 => (x"c1",x"02",x"6d",x"97"),
  1030 => (x"e8",x"c2",x"87",x"dc"),
  1031 => (x"74",x"49",x"bf",x"fc"),
  1032 => (x"de",x"fd",x"71",x"81"),
  1033 => (x"48",x"7e",x"70",x"87"),
  1034 => (x"f2",x"c0",x"02",x"98"),
  1035 => (x"c4",x"e9",x"c2",x"87"),
  1036 => (x"cb",x"4a",x"70",x"4b"),
  1037 => (x"ee",x"c1",x"ff",x"49"),
  1038 => (x"cb",x"4b",x"74",x"87"),
  1039 => (x"e7",x"e3",x"c1",x"93"),
  1040 => (x"c1",x"83",x"c4",x"83"),
  1041 => (x"74",x"7b",x"fa",x"c1"),
  1042 => (x"ef",x"c1",x"c1",x"49"),
  1043 => (x"c1",x"7b",x"75",x"87"),
  1044 => (x"bf",x"97",x"d4",x"e3"),
  1045 => (x"e9",x"c2",x"1e",x"49"),
  1046 => (x"e5",x"fd",x"49",x"c4"),
  1047 => (x"74",x"86",x"c4",x"87"),
  1048 => (x"d7",x"c1",x"c1",x"49"),
  1049 => (x"c1",x"49",x"c0",x"87"),
  1050 => (x"c2",x"87",x"f6",x"c2"),
  1051 => (x"c0",x"48",x"e4",x"e8"),
  1052 => (x"de",x"49",x"c1",x"78"),
  1053 => (x"fc",x"26",x"87",x"ca"),
  1054 => (x"6f",x"4c",x"87",x"c1"),
  1055 => (x"6e",x"69",x"64",x"61"),
  1056 => (x"2e",x"2e",x"2e",x"67"),
  1057 => (x"1e",x"73",x"1e",x"00"),
  1058 => (x"c2",x"49",x"4a",x"71"),
  1059 => (x"81",x"bf",x"fc",x"e8"),
  1060 => (x"87",x"ef",x"fb",x"71"),
  1061 => (x"02",x"9b",x"4b",x"70"),
  1062 => (x"e7",x"49",x"87",x"c4"),
  1063 => (x"e8",x"c2",x"87",x"e9"),
  1064 => (x"78",x"c0",x"48",x"fc"),
  1065 => (x"d7",x"dd",x"49",x"c1"),
  1066 => (x"87",x"d3",x"fb",x"87"),
  1067 => (x"c1",x"49",x"c0",x"1e"),
  1068 => (x"26",x"87",x"ee",x"c1"),
  1069 => (x"4a",x"71",x"1e",x"4f"),
  1070 => (x"c1",x"91",x"cb",x"49"),
  1071 => (x"c8",x"81",x"e7",x"e3"),
  1072 => (x"c2",x"48",x"11",x"81"),
  1073 => (x"c2",x"58",x"e8",x"e8"),
  1074 => (x"c0",x"48",x"fc",x"e8"),
  1075 => (x"dc",x"49",x"c1",x"78"),
  1076 => (x"4f",x"26",x"87",x"ee"),
  1077 => (x"02",x"99",x"71",x"1e"),
  1078 => (x"e4",x"c1",x"87",x"d2"),
  1079 => (x"50",x"c0",x"48",x"fc"),
  1080 => (x"c2",x"c1",x"80",x"f7"),
  1081 => (x"e3",x"c1",x"40",x"f5"),
  1082 => (x"87",x"ce",x"78",x"e0"),
  1083 => (x"48",x"f8",x"e4",x"c1"),
  1084 => (x"78",x"d9",x"e3",x"c1"),
  1085 => (x"c2",x"c1",x"80",x"fc"),
  1086 => (x"4f",x"26",x"78",x"ec"),
  1087 => (x"5c",x"5b",x"5e",x"0e"),
  1088 => (x"86",x"f4",x"0e",x"5d"),
  1089 => (x"4d",x"f2",x"db",x"c2"),
  1090 => (x"a6",x"c4",x"4c",x"c0"),
  1091 => (x"c2",x"78",x"c0",x"48"),
  1092 => (x"48",x"bf",x"fc",x"e8"),
  1093 => (x"c1",x"06",x"a8",x"c0"),
  1094 => (x"db",x"c2",x"87",x"c0"),
  1095 => (x"02",x"98",x"48",x"f2"),
  1096 => (x"c0",x"87",x"f7",x"c0"),
  1097 => (x"c8",x"1e",x"cf",x"f6"),
  1098 => (x"87",x"c7",x"02",x"66"),
  1099 => (x"c0",x"48",x"a6",x"c4"),
  1100 => (x"c4",x"87",x"c5",x"78"),
  1101 => (x"78",x"c1",x"48",x"a6"),
  1102 => (x"e6",x"49",x"66",x"c4"),
  1103 => (x"86",x"c4",x"87",x"c0"),
  1104 => (x"84",x"c1",x"4d",x"70"),
  1105 => (x"c1",x"48",x"66",x"c4"),
  1106 => (x"58",x"a6",x"c8",x"80"),
  1107 => (x"bf",x"fc",x"e8",x"c2"),
  1108 => (x"87",x"c6",x"03",x"ac"),
  1109 => (x"ff",x"05",x"9d",x"75"),
  1110 => (x"4c",x"c0",x"87",x"c9"),
  1111 => (x"c3",x"02",x"9d",x"75"),
  1112 => (x"f6",x"c0",x"87",x"dc"),
  1113 => (x"66",x"c8",x"1e",x"cf"),
  1114 => (x"cc",x"87",x"c7",x"02"),
  1115 => (x"78",x"c0",x"48",x"a6"),
  1116 => (x"a6",x"cc",x"87",x"c5"),
  1117 => (x"cc",x"78",x"c1",x"48"),
  1118 => (x"c1",x"e5",x"49",x"66"),
  1119 => (x"70",x"86",x"c4",x"87"),
  1120 => (x"02",x"98",x"48",x"7e"),
  1121 => (x"49",x"87",x"e4",x"c2"),
  1122 => (x"69",x"97",x"81",x"cb"),
  1123 => (x"02",x"99",x"d0",x"49"),
  1124 => (x"74",x"87",x"d4",x"c1"),
  1125 => (x"c1",x"91",x"cb",x"49"),
  1126 => (x"c1",x"81",x"e7",x"e3"),
  1127 => (x"c8",x"79",x"c5",x"c2"),
  1128 => (x"51",x"ff",x"c3",x"81"),
  1129 => (x"91",x"de",x"49",x"74"),
  1130 => (x"4d",x"d0",x"e9",x"c2"),
  1131 => (x"c1",x"c2",x"85",x"71"),
  1132 => (x"a5",x"c1",x"7d",x"97"),
  1133 => (x"51",x"e0",x"c0",x"49"),
  1134 => (x"97",x"c2",x"e4",x"c2"),
  1135 => (x"87",x"d2",x"02",x"bf"),
  1136 => (x"a5",x"c2",x"84",x"c1"),
  1137 => (x"c2",x"e4",x"c2",x"4b"),
  1138 => (x"fe",x"49",x"db",x"4a"),
  1139 => (x"c1",x"87",x"d8",x"fb"),
  1140 => (x"a5",x"cd",x"87",x"d9"),
  1141 => (x"c1",x"51",x"c0",x"49"),
  1142 => (x"4b",x"a5",x"c2",x"84"),
  1143 => (x"49",x"cb",x"4a",x"6e"),
  1144 => (x"87",x"c3",x"fb",x"fe"),
  1145 => (x"74",x"87",x"c4",x"c1"),
  1146 => (x"c1",x"91",x"cb",x"49"),
  1147 => (x"c1",x"81",x"e7",x"e3"),
  1148 => (x"c2",x"79",x"c2",x"c0"),
  1149 => (x"bf",x"97",x"c2",x"e4"),
  1150 => (x"74",x"87",x"d8",x"02"),
  1151 => (x"c1",x"91",x"de",x"49"),
  1152 => (x"d0",x"e9",x"c2",x"84"),
  1153 => (x"c2",x"83",x"71",x"4b"),
  1154 => (x"dd",x"4a",x"c2",x"e4"),
  1155 => (x"d6",x"fa",x"fe",x"49"),
  1156 => (x"74",x"87",x"d8",x"87"),
  1157 => (x"c2",x"93",x"de",x"4b"),
  1158 => (x"cb",x"83",x"d0",x"e9"),
  1159 => (x"51",x"c0",x"49",x"a3"),
  1160 => (x"6e",x"73",x"84",x"c1"),
  1161 => (x"fe",x"49",x"cb",x"4a"),
  1162 => (x"c4",x"87",x"fc",x"f9"),
  1163 => (x"80",x"c1",x"48",x"66"),
  1164 => (x"c7",x"58",x"a6",x"c8"),
  1165 => (x"c5",x"c0",x"03",x"ac"),
  1166 => (x"fc",x"05",x"6e",x"87"),
  1167 => (x"48",x"74",x"87",x"e4"),
  1168 => (x"f6",x"f4",x"8e",x"f4"),
  1169 => (x"1e",x"73",x"1e",x"87"),
  1170 => (x"cb",x"49",x"4b",x"71"),
  1171 => (x"e7",x"e3",x"c1",x"91"),
  1172 => (x"4a",x"a1",x"c8",x"81"),
  1173 => (x"48",x"d3",x"e3",x"c1"),
  1174 => (x"a1",x"c9",x"50",x"12"),
  1175 => (x"ee",x"f8",x"c0",x"4a"),
  1176 => (x"ca",x"50",x"12",x"48"),
  1177 => (x"d4",x"e3",x"c1",x"81"),
  1178 => (x"c1",x"50",x"11",x"48"),
  1179 => (x"bf",x"97",x"d4",x"e3"),
  1180 => (x"49",x"c0",x"1e",x"49"),
  1181 => (x"c2",x"87",x"cb",x"f5"),
  1182 => (x"de",x"48",x"e4",x"e8"),
  1183 => (x"d5",x"49",x"c1",x"78"),
  1184 => (x"f3",x"26",x"87",x"fe"),
  1185 => (x"5e",x"0e",x"87",x"f9"),
  1186 => (x"0e",x"5d",x"5c",x"5b"),
  1187 => (x"4d",x"71",x"86",x"f4"),
  1188 => (x"c1",x"91",x"cb",x"49"),
  1189 => (x"c8",x"81",x"e7",x"e3"),
  1190 => (x"a1",x"ca",x"4a",x"a1"),
  1191 => (x"48",x"a6",x"c4",x"7e"),
  1192 => (x"bf",x"ec",x"ec",x"c2"),
  1193 => (x"bf",x"97",x"6e",x"78"),
  1194 => (x"4c",x"66",x"c4",x"4b"),
  1195 => (x"48",x"12",x"2c",x"73"),
  1196 => (x"70",x"58",x"a6",x"cc"),
  1197 => (x"c9",x"84",x"c1",x"9c"),
  1198 => (x"49",x"69",x"97",x"81"),
  1199 => (x"c2",x"04",x"ac",x"b7"),
  1200 => (x"6e",x"4c",x"c0",x"87"),
  1201 => (x"c8",x"4a",x"bf",x"97"),
  1202 => (x"31",x"72",x"49",x"66"),
  1203 => (x"66",x"c4",x"b9",x"ff"),
  1204 => (x"72",x"48",x"74",x"99"),
  1205 => (x"48",x"4a",x"70",x"30"),
  1206 => (x"ec",x"c2",x"b0",x"71"),
  1207 => (x"e5",x"c0",x"58",x"f0"),
  1208 => (x"49",x"c0",x"87",x"da"),
  1209 => (x"75",x"87",x"d9",x"d4"),
  1210 => (x"cf",x"f7",x"c0",x"49"),
  1211 => (x"f2",x"8e",x"f4",x"87"),
  1212 => (x"73",x"1e",x"87",x"c9"),
  1213 => (x"49",x"4b",x"71",x"1e"),
  1214 => (x"73",x"87",x"cb",x"fe"),
  1215 => (x"87",x"c6",x"fe",x"49"),
  1216 => (x"1e",x"87",x"fc",x"f1"),
  1217 => (x"4b",x"71",x"1e",x"73"),
  1218 => (x"02",x"4a",x"a3",x"c6"),
  1219 => (x"c1",x"87",x"e3",x"c0"),
  1220 => (x"87",x"d6",x"02",x"8a"),
  1221 => (x"e8",x"c1",x"02",x"8a"),
  1222 => (x"c1",x"02",x"8a",x"87"),
  1223 => (x"02",x"8a",x"87",x"ca"),
  1224 => (x"8a",x"87",x"ef",x"c0"),
  1225 => (x"c1",x"87",x"d9",x"02"),
  1226 => (x"49",x"c7",x"87",x"e9"),
  1227 => (x"c1",x"87",x"c6",x"f6"),
  1228 => (x"e8",x"c2",x"87",x"ec"),
  1229 => (x"78",x"df",x"48",x"e4"),
  1230 => (x"c3",x"d3",x"49",x"c1"),
  1231 => (x"87",x"de",x"c1",x"87"),
  1232 => (x"bf",x"fc",x"e8",x"c2"),
  1233 => (x"87",x"cb",x"c1",x"02"),
  1234 => (x"c2",x"88",x"c1",x"48"),
  1235 => (x"c1",x"58",x"c0",x"e9"),
  1236 => (x"e9",x"c2",x"87",x"c1"),
  1237 => (x"c0",x"02",x"bf",x"c0"),
  1238 => (x"e8",x"c2",x"87",x"f9"),
  1239 => (x"c1",x"48",x"bf",x"fc"),
  1240 => (x"c0",x"e9",x"c2",x"80"),
  1241 => (x"87",x"eb",x"c0",x"58"),
  1242 => (x"bf",x"fc",x"e8",x"c2"),
  1243 => (x"c2",x"89",x"c6",x"49"),
  1244 => (x"c0",x"59",x"c0",x"e9"),
  1245 => (x"da",x"03",x"a9",x"b7"),
  1246 => (x"fc",x"e8",x"c2",x"87"),
  1247 => (x"d2",x"78",x"c0",x"48"),
  1248 => (x"c0",x"e9",x"c2",x"87"),
  1249 => (x"87",x"cb",x"02",x"bf"),
  1250 => (x"bf",x"fc",x"e8",x"c2"),
  1251 => (x"c2",x"80",x"c6",x"48"),
  1252 => (x"c0",x"58",x"c0",x"e9"),
  1253 => (x"87",x"e8",x"d1",x"49"),
  1254 => (x"f4",x"c0",x"49",x"73"),
  1255 => (x"de",x"ef",x"87",x"de"),
  1256 => (x"5b",x"5e",x"0e",x"87"),
  1257 => (x"ff",x"0e",x"5d",x"5c"),
  1258 => (x"a6",x"dc",x"86",x"d4"),
  1259 => (x"48",x"a6",x"c8",x"59"),
  1260 => (x"80",x"c4",x"78",x"c0"),
  1261 => (x"78",x"66",x"c0",x"c1"),
  1262 => (x"78",x"c1",x"80",x"c4"),
  1263 => (x"78",x"c1",x"80",x"c4"),
  1264 => (x"48",x"c0",x"e9",x"c2"),
  1265 => (x"e8",x"c2",x"78",x"c1"),
  1266 => (x"de",x"48",x"bf",x"e4"),
  1267 => (x"87",x"c9",x"05",x"a8"),
  1268 => (x"cc",x"87",x"e9",x"f4"),
  1269 => (x"e6",x"cf",x"58",x"a6"),
  1270 => (x"87",x"e2",x"e3",x"87"),
  1271 => (x"e3",x"87",x"c4",x"e4"),
  1272 => (x"4c",x"70",x"87",x"d1"),
  1273 => (x"02",x"ac",x"fb",x"c0"),
  1274 => (x"d8",x"87",x"fb",x"c1"),
  1275 => (x"ed",x"c1",x"05",x"66"),
  1276 => (x"66",x"fc",x"c0",x"87"),
  1277 => (x"6a",x"82",x"c4",x"4a"),
  1278 => (x"c1",x"1e",x"72",x"7e"),
  1279 => (x"c4",x"48",x"f4",x"df"),
  1280 => (x"a1",x"c8",x"49",x"66"),
  1281 => (x"71",x"41",x"20",x"4a"),
  1282 => (x"87",x"f9",x"05",x"aa"),
  1283 => (x"4a",x"26",x"51",x"10"),
  1284 => (x"48",x"66",x"fc",x"c0"),
  1285 => (x"78",x"c5",x"c9",x"c1"),
  1286 => (x"81",x"c7",x"49",x"6a"),
  1287 => (x"fc",x"c0",x"51",x"74"),
  1288 => (x"81",x"c8",x"49",x"66"),
  1289 => (x"fc",x"c0",x"51",x"c1"),
  1290 => (x"81",x"c9",x"49",x"66"),
  1291 => (x"fc",x"c0",x"51",x"c0"),
  1292 => (x"81",x"ca",x"49",x"66"),
  1293 => (x"1e",x"c1",x"51",x"c0"),
  1294 => (x"49",x"6a",x"1e",x"d8"),
  1295 => (x"f6",x"e2",x"81",x"c8"),
  1296 => (x"c1",x"86",x"c8",x"87"),
  1297 => (x"c0",x"48",x"66",x"c0"),
  1298 => (x"87",x"c7",x"01",x"a8"),
  1299 => (x"c1",x"48",x"a6",x"c8"),
  1300 => (x"c1",x"87",x"ce",x"78"),
  1301 => (x"c1",x"48",x"66",x"c0"),
  1302 => (x"58",x"a6",x"d0",x"88"),
  1303 => (x"c2",x"e2",x"87",x"c3"),
  1304 => (x"48",x"a6",x"d0",x"87"),
  1305 => (x"9c",x"74",x"78",x"c2"),
  1306 => (x"87",x"cf",x"cd",x"02"),
  1307 => (x"c1",x"48",x"66",x"c8"),
  1308 => (x"03",x"a8",x"66",x"c4"),
  1309 => (x"dc",x"87",x"c4",x"cd"),
  1310 => (x"78",x"c0",x"48",x"a6"),
  1311 => (x"78",x"c0",x"80",x"e8"),
  1312 => (x"70",x"87",x"f0",x"e0"),
  1313 => (x"ac",x"d0",x"c1",x"4c"),
  1314 => (x"87",x"d7",x"c2",x"05"),
  1315 => (x"e3",x"7e",x"66",x"c4"),
  1316 => (x"a6",x"c8",x"87",x"d4"),
  1317 => (x"87",x"db",x"e0",x"58"),
  1318 => (x"ec",x"c0",x"4c",x"70"),
  1319 => (x"ed",x"c1",x"05",x"ac"),
  1320 => (x"49",x"66",x"c8",x"87"),
  1321 => (x"fc",x"c0",x"91",x"cb"),
  1322 => (x"a1",x"c4",x"81",x"66"),
  1323 => (x"c8",x"4d",x"6a",x"4a"),
  1324 => (x"66",x"c4",x"4a",x"a1"),
  1325 => (x"f5",x"c2",x"c1",x"52"),
  1326 => (x"f6",x"df",x"ff",x"79"),
  1327 => (x"9c",x"4c",x"70",x"87"),
  1328 => (x"c0",x"87",x"d9",x"02"),
  1329 => (x"d3",x"02",x"ac",x"fb"),
  1330 => (x"ff",x"55",x"74",x"87"),
  1331 => (x"70",x"87",x"e4",x"df"),
  1332 => (x"c7",x"02",x"9c",x"4c"),
  1333 => (x"ac",x"fb",x"c0",x"87"),
  1334 => (x"87",x"ed",x"ff",x"05"),
  1335 => (x"c2",x"55",x"e0",x"c0"),
  1336 => (x"97",x"c0",x"55",x"c1"),
  1337 => (x"48",x"66",x"d8",x"7d"),
  1338 => (x"db",x"05",x"a8",x"6e"),
  1339 => (x"48",x"66",x"c8",x"87"),
  1340 => (x"04",x"a8",x"66",x"cc"),
  1341 => (x"66",x"c8",x"87",x"ca"),
  1342 => (x"cc",x"80",x"c1",x"48"),
  1343 => (x"87",x"c8",x"58",x"a6"),
  1344 => (x"c1",x"48",x"66",x"cc"),
  1345 => (x"58",x"a6",x"d0",x"88"),
  1346 => (x"87",x"e7",x"de",x"ff"),
  1347 => (x"d0",x"c1",x"4c",x"70"),
  1348 => (x"87",x"c8",x"05",x"ac"),
  1349 => (x"c1",x"48",x"66",x"d4"),
  1350 => (x"58",x"a6",x"d8",x"80"),
  1351 => (x"02",x"ac",x"d0",x"c1"),
  1352 => (x"c4",x"87",x"e9",x"fd"),
  1353 => (x"66",x"d8",x"48",x"66"),
  1354 => (x"e0",x"c9",x"05",x"a8"),
  1355 => (x"a6",x"e0",x"c0",x"87"),
  1356 => (x"74",x"78",x"c0",x"48"),
  1357 => (x"88",x"fb",x"c0",x"48"),
  1358 => (x"98",x"48",x"7e",x"70"),
  1359 => (x"87",x"e2",x"c9",x"02"),
  1360 => (x"70",x"88",x"cb",x"48"),
  1361 => (x"02",x"98",x"48",x"7e"),
  1362 => (x"48",x"87",x"cd",x"c1"),
  1363 => (x"7e",x"70",x"88",x"c9"),
  1364 => (x"c3",x"02",x"98",x"48"),
  1365 => (x"c4",x"48",x"87",x"fe"),
  1366 => (x"48",x"7e",x"70",x"88"),
  1367 => (x"87",x"ce",x"02",x"98"),
  1368 => (x"70",x"88",x"c1",x"48"),
  1369 => (x"02",x"98",x"48",x"7e"),
  1370 => (x"c8",x"87",x"e9",x"c3"),
  1371 => (x"a6",x"dc",x"87",x"d6"),
  1372 => (x"78",x"f0",x"c0",x"48"),
  1373 => (x"87",x"fb",x"dc",x"ff"),
  1374 => (x"ec",x"c0",x"4c",x"70"),
  1375 => (x"c4",x"c0",x"02",x"ac"),
  1376 => (x"a6",x"e0",x"c0",x"87"),
  1377 => (x"ac",x"ec",x"c0",x"5c"),
  1378 => (x"ff",x"87",x"cd",x"02"),
  1379 => (x"70",x"87",x"e4",x"dc"),
  1380 => (x"ac",x"ec",x"c0",x"4c"),
  1381 => (x"87",x"f3",x"ff",x"05"),
  1382 => (x"02",x"ac",x"ec",x"c0"),
  1383 => (x"ff",x"87",x"c4",x"c0"),
  1384 => (x"c0",x"87",x"d0",x"dc"),
  1385 => (x"d0",x"1e",x"ca",x"1e"),
  1386 => (x"91",x"cb",x"49",x"66"),
  1387 => (x"48",x"66",x"c4",x"c1"),
  1388 => (x"a6",x"cc",x"80",x"71"),
  1389 => (x"48",x"66",x"c8",x"58"),
  1390 => (x"a6",x"d0",x"80",x"c4"),
  1391 => (x"bf",x"66",x"cc",x"58"),
  1392 => (x"f2",x"dc",x"ff",x"49"),
  1393 => (x"de",x"1e",x"c1",x"87"),
  1394 => (x"bf",x"66",x"d4",x"1e"),
  1395 => (x"e6",x"dc",x"ff",x"49"),
  1396 => (x"70",x"86",x"d0",x"87"),
  1397 => (x"08",x"c0",x"48",x"49"),
  1398 => (x"a6",x"e8",x"c0",x"88"),
  1399 => (x"06",x"a8",x"c0",x"58"),
  1400 => (x"c0",x"87",x"ee",x"c0"),
  1401 => (x"dd",x"48",x"66",x"e4"),
  1402 => (x"e4",x"c0",x"03",x"a8"),
  1403 => (x"bf",x"66",x"c4",x"87"),
  1404 => (x"66",x"e4",x"c0",x"49"),
  1405 => (x"51",x"e0",x"c0",x"81"),
  1406 => (x"49",x"66",x"e4",x"c0"),
  1407 => (x"66",x"c4",x"81",x"c1"),
  1408 => (x"c1",x"c2",x"81",x"bf"),
  1409 => (x"66",x"e4",x"c0",x"51"),
  1410 => (x"c4",x"81",x"c2",x"49"),
  1411 => (x"c0",x"81",x"bf",x"66"),
  1412 => (x"c1",x"48",x"6e",x"51"),
  1413 => (x"6e",x"78",x"c5",x"c9"),
  1414 => (x"d0",x"81",x"c8",x"49"),
  1415 => (x"49",x"6e",x"51",x"66"),
  1416 => (x"66",x"d4",x"81",x"c9"),
  1417 => (x"ca",x"49",x"6e",x"51"),
  1418 => (x"51",x"66",x"dc",x"81"),
  1419 => (x"c1",x"48",x"66",x"d0"),
  1420 => (x"58",x"a6",x"d4",x"80"),
  1421 => (x"cc",x"48",x"66",x"c8"),
  1422 => (x"c0",x"04",x"a8",x"66"),
  1423 => (x"66",x"c8",x"87",x"cb"),
  1424 => (x"cc",x"80",x"c1",x"48"),
  1425 => (x"d9",x"c5",x"58",x"a6"),
  1426 => (x"48",x"66",x"cc",x"87"),
  1427 => (x"a6",x"d0",x"88",x"c1"),
  1428 => (x"87",x"ce",x"c5",x"58"),
  1429 => (x"87",x"ce",x"dc",x"ff"),
  1430 => (x"58",x"a6",x"e8",x"c0"),
  1431 => (x"87",x"c6",x"dc",x"ff"),
  1432 => (x"58",x"a6",x"e0",x"c0"),
  1433 => (x"05",x"a8",x"ec",x"c0"),
  1434 => (x"dc",x"87",x"ca",x"c0"),
  1435 => (x"e4",x"c0",x"48",x"a6"),
  1436 => (x"c4",x"c0",x"78",x"66"),
  1437 => (x"fa",x"d8",x"ff",x"87"),
  1438 => (x"49",x"66",x"c8",x"87"),
  1439 => (x"fc",x"c0",x"91",x"cb"),
  1440 => (x"80",x"71",x"48",x"66"),
  1441 => (x"c8",x"4a",x"7e",x"70"),
  1442 => (x"ca",x"49",x"6e",x"82"),
  1443 => (x"66",x"e4",x"c0",x"81"),
  1444 => (x"49",x"66",x"dc",x"51"),
  1445 => (x"e4",x"c0",x"81",x"c1"),
  1446 => (x"48",x"c1",x"89",x"66"),
  1447 => (x"49",x"70",x"30",x"71"),
  1448 => (x"97",x"71",x"89",x"c1"),
  1449 => (x"ec",x"ec",x"c2",x"7a"),
  1450 => (x"e4",x"c0",x"49",x"bf"),
  1451 => (x"6a",x"97",x"29",x"66"),
  1452 => (x"98",x"71",x"48",x"4a"),
  1453 => (x"58",x"a6",x"ec",x"c0"),
  1454 => (x"81",x"c4",x"49",x"6e"),
  1455 => (x"66",x"d8",x"4d",x"69"),
  1456 => (x"a8",x"66",x"c4",x"48"),
  1457 => (x"87",x"c8",x"c0",x"02"),
  1458 => (x"c0",x"48",x"a6",x"c4"),
  1459 => (x"87",x"c5",x"c0",x"78"),
  1460 => (x"c1",x"48",x"a6",x"c4"),
  1461 => (x"1e",x"66",x"c4",x"78"),
  1462 => (x"75",x"1e",x"e0",x"c0"),
  1463 => (x"d6",x"d8",x"ff",x"49"),
  1464 => (x"70",x"86",x"c8",x"87"),
  1465 => (x"ac",x"b7",x"c0",x"4c"),
  1466 => (x"87",x"d4",x"c1",x"06"),
  1467 => (x"e0",x"c0",x"85",x"74"),
  1468 => (x"75",x"89",x"74",x"49"),
  1469 => (x"fd",x"df",x"c1",x"4b"),
  1470 => (x"e6",x"fe",x"71",x"4a"),
  1471 => (x"85",x"c2",x"87",x"e9"),
  1472 => (x"48",x"66",x"e0",x"c0"),
  1473 => (x"e4",x"c0",x"80",x"c1"),
  1474 => (x"e8",x"c0",x"58",x"a6"),
  1475 => (x"81",x"c1",x"49",x"66"),
  1476 => (x"c0",x"02",x"a9",x"70"),
  1477 => (x"a6",x"c4",x"87",x"c8"),
  1478 => (x"c0",x"78",x"c0",x"48"),
  1479 => (x"a6",x"c4",x"87",x"c5"),
  1480 => (x"c4",x"78",x"c1",x"48"),
  1481 => (x"a4",x"c2",x"1e",x"66"),
  1482 => (x"48",x"e0",x"c0",x"49"),
  1483 => (x"49",x"70",x"88",x"71"),
  1484 => (x"ff",x"49",x"75",x"1e"),
  1485 => (x"c8",x"87",x"c0",x"d7"),
  1486 => (x"a8",x"b7",x"c0",x"86"),
  1487 => (x"87",x"c0",x"ff",x"01"),
  1488 => (x"02",x"66",x"e0",x"c0"),
  1489 => (x"6e",x"87",x"d1",x"c0"),
  1490 => (x"c0",x"81",x"c9",x"49"),
  1491 => (x"6e",x"51",x"66",x"e0"),
  1492 => (x"c6",x"ca",x"c1",x"48"),
  1493 => (x"87",x"cc",x"c0",x"78"),
  1494 => (x"81",x"c9",x"49",x"6e"),
  1495 => (x"48",x"6e",x"51",x"c2"),
  1496 => (x"78",x"f2",x"cb",x"c1"),
  1497 => (x"cc",x"48",x"66",x"c8"),
  1498 => (x"c0",x"04",x"a8",x"66"),
  1499 => (x"66",x"c8",x"87",x"cb"),
  1500 => (x"cc",x"80",x"c1",x"48"),
  1501 => (x"e9",x"c0",x"58",x"a6"),
  1502 => (x"48",x"66",x"cc",x"87"),
  1503 => (x"a6",x"d0",x"88",x"c1"),
  1504 => (x"87",x"de",x"c0",x"58"),
  1505 => (x"87",x"db",x"d5",x"ff"),
  1506 => (x"d5",x"c0",x"4c",x"70"),
  1507 => (x"ac",x"c6",x"c1",x"87"),
  1508 => (x"87",x"c8",x"c0",x"05"),
  1509 => (x"c1",x"48",x"66",x"d0"),
  1510 => (x"58",x"a6",x"d4",x"80"),
  1511 => (x"87",x"c3",x"d5",x"ff"),
  1512 => (x"66",x"d4",x"4c",x"70"),
  1513 => (x"d8",x"80",x"c1",x"48"),
  1514 => (x"9c",x"74",x"58",x"a6"),
  1515 => (x"87",x"cb",x"c0",x"02"),
  1516 => (x"c1",x"48",x"66",x"c8"),
  1517 => (x"04",x"a8",x"66",x"c4"),
  1518 => (x"ff",x"87",x"fc",x"f2"),
  1519 => (x"c8",x"87",x"db",x"d4"),
  1520 => (x"a8",x"c7",x"48",x"66"),
  1521 => (x"87",x"e5",x"c0",x"03"),
  1522 => (x"48",x"c0",x"e9",x"c2"),
  1523 => (x"66",x"c8",x"78",x"c0"),
  1524 => (x"c0",x"91",x"cb",x"49"),
  1525 => (x"c4",x"81",x"66",x"fc"),
  1526 => (x"4a",x"6a",x"4a",x"a1"),
  1527 => (x"c8",x"79",x"52",x"c0"),
  1528 => (x"80",x"c1",x"48",x"66"),
  1529 => (x"c7",x"58",x"a6",x"cc"),
  1530 => (x"db",x"ff",x"04",x"a8"),
  1531 => (x"8e",x"d4",x"ff",x"87"),
  1532 => (x"87",x"c7",x"de",x"ff"),
  1533 => (x"64",x"61",x"6f",x"4c"),
  1534 => (x"20",x"2e",x"2a",x"20"),
  1535 => (x"00",x"20",x"3a",x"00"),
  1536 => (x"71",x"1e",x"73",x"1e"),
  1537 => (x"c6",x"02",x"9b",x"4b"),
  1538 => (x"fc",x"e8",x"c2",x"87"),
  1539 => (x"c7",x"78",x"c0",x"48"),
  1540 => (x"fc",x"e8",x"c2",x"1e"),
  1541 => (x"e3",x"c1",x"1e",x"bf"),
  1542 => (x"e8",x"c2",x"1e",x"e7"),
  1543 => (x"ed",x"49",x"bf",x"e4"),
  1544 => (x"86",x"cc",x"87",x"ff"),
  1545 => (x"bf",x"e4",x"e8",x"c2"),
  1546 => (x"87",x"e8",x"e2",x"49"),
  1547 => (x"c8",x"02",x"9b",x"73"),
  1548 => (x"e7",x"e3",x"c1",x"87"),
  1549 => (x"d5",x"e3",x"c0",x"49"),
  1550 => (x"c2",x"dd",x"ff",x"87"),
  1551 => (x"e3",x"c1",x"1e",x"87"),
  1552 => (x"50",x"c0",x"48",x"d3"),
  1553 => (x"bf",x"ca",x"e5",x"c1"),
  1554 => (x"e2",x"d7",x"ff",x"49"),
  1555 => (x"26",x"48",x"c0",x"87"),
  1556 => (x"d9",x"c7",x"1e",x"4f"),
  1557 => (x"fe",x"49",x"c1",x"87"),
  1558 => (x"e9",x"c2",x"87",x"e6"),
  1559 => (x"50",x"c0",x"48",x"c4"),
  1560 => (x"87",x"f3",x"e9",x"fe"),
  1561 => (x"cd",x"02",x"98",x"70"),
  1562 => (x"ed",x"f2",x"fe",x"87"),
  1563 => (x"02",x"98",x"70",x"87"),
  1564 => (x"4a",x"c1",x"87",x"c4"),
  1565 => (x"4a",x"c0",x"87",x"c2"),
  1566 => (x"ce",x"05",x"9a",x"72"),
  1567 => (x"c1",x"1e",x"c0",x"87"),
  1568 => (x"c0",x"49",x"fd",x"e2"),
  1569 => (x"c4",x"87",x"fb",x"ef"),
  1570 => (x"c2",x"87",x"fe",x"86"),
  1571 => (x"c0",x"48",x"fc",x"e8"),
  1572 => (x"e4",x"e8",x"c2",x"78"),
  1573 => (x"1e",x"78",x"c0",x"48"),
  1574 => (x"49",x"c8",x"e3",x"c1"),
  1575 => (x"87",x"e2",x"ef",x"c0"),
  1576 => (x"d8",x"fe",x"1e",x"c0"),
  1577 => (x"c0",x"49",x"70",x"87"),
  1578 => (x"c8",x"87",x"d7",x"ef"),
  1579 => (x"87",x"fd",x"c2",x"86"),
  1580 => (x"87",x"d7",x"e3",x"c0"),
  1581 => (x"87",x"c4",x"f3",x"c0"),
  1582 => (x"26",x"87",x"f5",x"ff"),
  1583 => (x"20",x"44",x"53",x"4f"),
  1584 => (x"6c",x"69",x"61",x"66"),
  1585 => (x"00",x"2e",x"64",x"65"),
  1586 => (x"74",x"6f",x"6f",x"42"),
  1587 => (x"2e",x"67",x"6e",x"69"),
  1588 => (x"00",x"00",x"2e",x"2e"),
  1589 => (x"00",x"00",x"01",x"00"),
  1590 => (x"45",x"20",x"80",x"00"),
  1591 => (x"00",x"74",x"69",x"78"),
  1592 => (x"61",x"42",x"20",x"80"),
  1593 => (x"02",x"00",x"6b",x"63"),
  1594 => (x"50",x"00",x"00",x"10"),
  1595 => (x"00",x"00",x"00",x"2a"),
  1596 => (x"10",x"02",x"00",x"00"),
  1597 => (x"2a",x"6e",x"00",x"00"),
  1598 => (x"00",x"00",x"00",x"00"),
  1599 => (x"00",x"10",x"02",x"00"),
  1600 => (x"00",x"2a",x"8c",x"00"),
  1601 => (x"00",x"00",x"00",x"00"),
  1602 => (x"00",x"00",x"10",x"02"),
  1603 => (x"00",x"00",x"2a",x"aa"),
  1604 => (x"02",x"00",x"00",x"00"),
  1605 => (x"c8",x"00",x"00",x"10"),
  1606 => (x"00",x"00",x"00",x"2a"),
  1607 => (x"10",x"02",x"00",x"00"),
  1608 => (x"2a",x"e6",x"00",x"00"),
  1609 => (x"00",x"00",x"00",x"00"),
  1610 => (x"00",x"10",x"02",x"00"),
  1611 => (x"00",x"2b",x"04",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"00",x"10",x"b5"),
  1614 => (x"00",x"00",x"00",x"00"),
  1615 => (x"03",x"00",x"00",x"00"),
  1616 => (x"00",x"00",x"00",x"13"),
  1617 => (x"00",x"00",x"00",x"00"),
  1618 => (x"19",x"4e",x"00",x"00"),
  1619 => (x"4f",x"42",x"00",x"00"),
  1620 => (x"20",x"20",x"54",x"4f"),
  1621 => (x"4f",x"52",x"20",x"20"),
  1622 => (x"fe",x"1e",x"00",x"4d"),
  1623 => (x"78",x"c0",x"48",x"f0"),
  1624 => (x"09",x"79",x"09",x"cd"),
  1625 => (x"fe",x"1e",x"4f",x"26"),
  1626 => (x"26",x"48",x"bf",x"f0"),
  1627 => (x"f0",x"fe",x"1e",x"4f"),
  1628 => (x"26",x"78",x"c1",x"48"),
  1629 => (x"f0",x"fe",x"1e",x"4f"),
  1630 => (x"26",x"78",x"c0",x"48"),
  1631 => (x"4a",x"71",x"1e",x"4f"),
  1632 => (x"26",x"51",x"52",x"c0"),
  1633 => (x"5b",x"5e",x"0e",x"4f"),
  1634 => (x"f4",x"0e",x"5d",x"5c"),
  1635 => (x"97",x"4d",x"71",x"86"),
  1636 => (x"a5",x"c1",x"7e",x"6d"),
  1637 => (x"48",x"6c",x"97",x"4c"),
  1638 => (x"6e",x"58",x"a6",x"c8"),
  1639 => (x"a8",x"66",x"c4",x"48"),
  1640 => (x"ff",x"87",x"c5",x"05"),
  1641 => (x"87",x"e6",x"c0",x"48"),
  1642 => (x"c2",x"87",x"ca",x"ff"),
  1643 => (x"6c",x"97",x"49",x"a5"),
  1644 => (x"4b",x"a3",x"71",x"4b"),
  1645 => (x"97",x"4b",x"6b",x"97"),
  1646 => (x"48",x"6e",x"7e",x"6c"),
  1647 => (x"a6",x"c8",x"80",x"c1"),
  1648 => (x"cc",x"98",x"c7",x"58"),
  1649 => (x"97",x"70",x"58",x"a6"),
  1650 => (x"87",x"e1",x"fe",x"7c"),
  1651 => (x"8e",x"f4",x"48",x"73"),
  1652 => (x"4c",x"26",x"4d",x"26"),
  1653 => (x"4f",x"26",x"4b",x"26"),
  1654 => (x"5c",x"5b",x"5e",x"0e"),
  1655 => (x"71",x"86",x"f4",x"0e"),
  1656 => (x"4a",x"66",x"d8",x"4c"),
  1657 => (x"c2",x"9a",x"ff",x"c3"),
  1658 => (x"6c",x"97",x"4b",x"a4"),
  1659 => (x"49",x"a1",x"73",x"49"),
  1660 => (x"6c",x"97",x"51",x"72"),
  1661 => (x"c1",x"48",x"6e",x"7e"),
  1662 => (x"58",x"a6",x"c8",x"80"),
  1663 => (x"a6",x"cc",x"98",x"c7"),
  1664 => (x"f4",x"54",x"70",x"58"),
  1665 => (x"87",x"ca",x"ff",x"8e"),
  1666 => (x"e8",x"fd",x"1e",x"1e"),
  1667 => (x"4a",x"bf",x"e0",x"87"),
  1668 => (x"c0",x"e0",x"c0",x"49"),
  1669 => (x"87",x"cb",x"02",x"99"),
  1670 => (x"ec",x"c2",x"1e",x"72"),
  1671 => (x"f7",x"fe",x"49",x"e2"),
  1672 => (x"fd",x"86",x"c4",x"87"),
  1673 => (x"7e",x"70",x"87",x"c0"),
  1674 => (x"26",x"87",x"c2",x"fd"),
  1675 => (x"c2",x"1e",x"4f",x"26"),
  1676 => (x"fd",x"49",x"e2",x"ec"),
  1677 => (x"e8",x"c1",x"87",x"c7"),
  1678 => (x"dd",x"fc",x"49",x"c8"),
  1679 => (x"87",x"ee",x"c3",x"87"),
  1680 => (x"5e",x"0e",x"4f",x"26"),
  1681 => (x"0e",x"5d",x"5c",x"5b"),
  1682 => (x"ec",x"c2",x"4d",x"71"),
  1683 => (x"f4",x"fc",x"49",x"e2"),
  1684 => (x"c0",x"4b",x"70",x"87"),
  1685 => (x"c3",x"04",x"ab",x"b7"),
  1686 => (x"f0",x"c3",x"87",x"c2"),
  1687 => (x"87",x"c9",x"05",x"ab"),
  1688 => (x"48",x"e6",x"ec",x"c1"),
  1689 => (x"e3",x"c2",x"78",x"c1"),
  1690 => (x"ab",x"e0",x"c3",x"87"),
  1691 => (x"c1",x"87",x"c9",x"05"),
  1692 => (x"c1",x"48",x"ea",x"ec"),
  1693 => (x"87",x"d4",x"c2",x"78"),
  1694 => (x"bf",x"ea",x"ec",x"c1"),
  1695 => (x"c2",x"87",x"c6",x"02"),
  1696 => (x"c2",x"4c",x"a3",x"c0"),
  1697 => (x"c1",x"4c",x"73",x"87"),
  1698 => (x"02",x"bf",x"e6",x"ec"),
  1699 => (x"74",x"87",x"e0",x"c0"),
  1700 => (x"29",x"b7",x"c4",x"49"),
  1701 => (x"fd",x"ed",x"c1",x"91"),
  1702 => (x"cf",x"4a",x"74",x"81"),
  1703 => (x"c1",x"92",x"c2",x"9a"),
  1704 => (x"70",x"30",x"72",x"48"),
  1705 => (x"72",x"ba",x"ff",x"4a"),
  1706 => (x"70",x"98",x"69",x"48"),
  1707 => (x"74",x"87",x"db",x"79"),
  1708 => (x"29",x"b7",x"c4",x"49"),
  1709 => (x"fd",x"ed",x"c1",x"91"),
  1710 => (x"cf",x"4a",x"74",x"81"),
  1711 => (x"c3",x"92",x"c2",x"9a"),
  1712 => (x"70",x"30",x"72",x"48"),
  1713 => (x"b0",x"69",x"48",x"4a"),
  1714 => (x"9d",x"75",x"79",x"70"),
  1715 => (x"87",x"f0",x"c0",x"05"),
  1716 => (x"c8",x"48",x"d0",x"ff"),
  1717 => (x"d4",x"ff",x"78",x"e1"),
  1718 => (x"c1",x"78",x"c5",x"48"),
  1719 => (x"02",x"bf",x"ea",x"ec"),
  1720 => (x"e0",x"c3",x"87",x"c3"),
  1721 => (x"e6",x"ec",x"c1",x"78"),
  1722 => (x"87",x"c6",x"02",x"bf"),
  1723 => (x"c3",x"48",x"d4",x"ff"),
  1724 => (x"d4",x"ff",x"78",x"f0"),
  1725 => (x"ff",x"0b",x"7b",x"0b"),
  1726 => (x"e1",x"c8",x"48",x"d0"),
  1727 => (x"78",x"e0",x"c0",x"78"),
  1728 => (x"48",x"ea",x"ec",x"c1"),
  1729 => (x"ec",x"c1",x"78",x"c0"),
  1730 => (x"78",x"c0",x"48",x"e6"),
  1731 => (x"49",x"e2",x"ec",x"c2"),
  1732 => (x"70",x"87",x"f2",x"f9"),
  1733 => (x"ab",x"b7",x"c0",x"4b"),
  1734 => (x"87",x"fe",x"fc",x"03"),
  1735 => (x"4d",x"26",x"48",x"c0"),
  1736 => (x"4b",x"26",x"4c",x"26"),
  1737 => (x"00",x"00",x"4f",x"26"),
  1738 => (x"00",x"00",x"00",x"00"),
  1739 => (x"c0",x"1e",x"00",x"00"),
  1740 => (x"c4",x"49",x"72",x"4a"),
  1741 => (x"fd",x"ed",x"c1",x"91"),
  1742 => (x"c1",x"79",x"c0",x"81"),
  1743 => (x"aa",x"b7",x"d0",x"82"),
  1744 => (x"26",x"87",x"ee",x"04"),
  1745 => (x"5b",x"5e",x"0e",x"4f"),
  1746 => (x"71",x"0e",x"5d",x"5c"),
  1747 => (x"87",x"e5",x"f8",x"4d"),
  1748 => (x"b7",x"c4",x"4a",x"75"),
  1749 => (x"ed",x"c1",x"92",x"2a"),
  1750 => (x"4c",x"75",x"82",x"fd"),
  1751 => (x"94",x"c2",x"9c",x"cf"),
  1752 => (x"74",x"4b",x"49",x"6a"),
  1753 => (x"c2",x"9b",x"c3",x"2b"),
  1754 => (x"70",x"30",x"74",x"48"),
  1755 => (x"74",x"bc",x"ff",x"4c"),
  1756 => (x"70",x"98",x"71",x"48"),
  1757 => (x"87",x"f5",x"f7",x"7a"),
  1758 => (x"e1",x"fe",x"48",x"73"),
  1759 => (x"00",x"00",x"00",x"87"),
  1760 => (x"00",x"00",x"00",x"00"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"00",x"00"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"00",x"00",x"00",x"00"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"d0",x"ff",x"1e",x"00"),
  1776 => (x"78",x"e1",x"c8",x"48"),
  1777 => (x"d4",x"ff",x"48",x"71"),
  1778 => (x"4f",x"26",x"78",x"08"),
  1779 => (x"48",x"d0",x"ff",x"1e"),
  1780 => (x"71",x"78",x"e1",x"c8"),
  1781 => (x"08",x"d4",x"ff",x"48"),
  1782 => (x"48",x"66",x"c4",x"78"),
  1783 => (x"78",x"08",x"d4",x"ff"),
  1784 => (x"71",x"1e",x"4f",x"26"),
  1785 => (x"49",x"66",x"c4",x"4a"),
  1786 => (x"ff",x"49",x"72",x"1e"),
  1787 => (x"d0",x"ff",x"87",x"de"),
  1788 => (x"78",x"e0",x"c0",x"48"),
  1789 => (x"1e",x"4f",x"26",x"26"),
  1790 => (x"4b",x"71",x"1e",x"73"),
  1791 => (x"1e",x"49",x"66",x"c8"),
  1792 => (x"e0",x"c1",x"4a",x"73"),
  1793 => (x"d9",x"ff",x"49",x"a2"),
  1794 => (x"87",x"c4",x"26",x"87"),
  1795 => (x"4c",x"26",x"4d",x"26"),
  1796 => (x"4f",x"26",x"4b",x"26"),
  1797 => (x"71",x"1e",x"73",x"1e"),
  1798 => (x"b7",x"c2",x"4b",x"4a"),
  1799 => (x"87",x"c8",x"03",x"ab"),
  1800 => (x"c3",x"4a",x"49",x"a3"),
  1801 => (x"87",x"c7",x"9a",x"ff"),
  1802 => (x"4a",x"49",x"a3",x"ce"),
  1803 => (x"c8",x"9a",x"ff",x"c3"),
  1804 => (x"72",x"1e",x"49",x"66"),
  1805 => (x"87",x"ea",x"fe",x"49"),
  1806 => (x"87",x"d4",x"ff",x"26"),
  1807 => (x"4a",x"d4",x"ff",x"1e"),
  1808 => (x"ff",x"7a",x"ff",x"c3"),
  1809 => (x"e1",x"c0",x"48",x"d0"),
  1810 => (x"c2",x"7a",x"de",x"78"),
  1811 => (x"7a",x"bf",x"ec",x"ec"),
  1812 => (x"28",x"c8",x"48",x"49"),
  1813 => (x"48",x"71",x"7a",x"70"),
  1814 => (x"7a",x"70",x"28",x"d0"),
  1815 => (x"28",x"d8",x"48",x"71"),
  1816 => (x"d0",x"ff",x"7a",x"70"),
  1817 => (x"78",x"e0",x"c0",x"48"),
  1818 => (x"ff",x"1e",x"4f",x"26"),
  1819 => (x"c9",x"c8",x"48",x"d0"),
  1820 => (x"ff",x"48",x"71",x"78"),
  1821 => (x"26",x"78",x"08",x"d4"),
  1822 => (x"4a",x"71",x"1e",x"4f"),
  1823 => (x"ff",x"87",x"eb",x"49"),
  1824 => (x"78",x"c8",x"48",x"d0"),
  1825 => (x"73",x"1e",x"4f",x"26"),
  1826 => (x"c2",x"4b",x"71",x"1e"),
  1827 => (x"02",x"bf",x"fc",x"ec"),
  1828 => (x"eb",x"c2",x"87",x"c3"),
  1829 => (x"48",x"d0",x"ff",x"87"),
  1830 => (x"73",x"78",x"c9",x"c8"),
  1831 => (x"b0",x"e0",x"c0",x"48"),
  1832 => (x"78",x"08",x"d4",x"ff"),
  1833 => (x"48",x"f0",x"ec",x"c2"),
  1834 => (x"66",x"c8",x"78",x"c0"),
  1835 => (x"c3",x"87",x"c5",x"02"),
  1836 => (x"87",x"c2",x"49",x"ff"),
  1837 => (x"ec",x"c2",x"49",x"c0"),
  1838 => (x"66",x"cc",x"59",x"f8"),
  1839 => (x"c5",x"87",x"c6",x"02"),
  1840 => (x"c4",x"4a",x"d5",x"d5"),
  1841 => (x"ff",x"ff",x"cf",x"87"),
  1842 => (x"fc",x"ec",x"c2",x"4a"),
  1843 => (x"fc",x"ec",x"c2",x"5a"),
  1844 => (x"c4",x"78",x"c1",x"48"),
  1845 => (x"26",x"4d",x"26",x"87"),
  1846 => (x"26",x"4b",x"26",x"4c"),
  1847 => (x"5b",x"5e",x"0e",x"4f"),
  1848 => (x"71",x"0e",x"5d",x"5c"),
  1849 => (x"f8",x"ec",x"c2",x"4a"),
  1850 => (x"9a",x"72",x"4c",x"bf"),
  1851 => (x"49",x"87",x"cb",x"02"),
  1852 => (x"f1",x"c1",x"91",x"c8"),
  1853 => (x"83",x"71",x"4b",x"fc"),
  1854 => (x"f5",x"c1",x"87",x"c4"),
  1855 => (x"4d",x"c0",x"4b",x"fc"),
  1856 => (x"99",x"74",x"49",x"13"),
  1857 => (x"bf",x"f4",x"ec",x"c2"),
  1858 => (x"ff",x"b8",x"71",x"48"),
  1859 => (x"c1",x"78",x"08",x"d4"),
  1860 => (x"c8",x"85",x"2c",x"b7"),
  1861 => (x"e7",x"04",x"ad",x"b7"),
  1862 => (x"f0",x"ec",x"c2",x"87"),
  1863 => (x"80",x"c8",x"48",x"bf"),
  1864 => (x"58",x"f4",x"ec",x"c2"),
  1865 => (x"1e",x"87",x"ee",x"fe"),
  1866 => (x"4b",x"71",x"1e",x"73"),
  1867 => (x"02",x"9a",x"4a",x"13"),
  1868 => (x"49",x"72",x"87",x"cb"),
  1869 => (x"13",x"87",x"e6",x"fe"),
  1870 => (x"f5",x"05",x"9a",x"4a"),
  1871 => (x"87",x"d9",x"fe",x"87"),
  1872 => (x"f0",x"ec",x"c2",x"1e"),
  1873 => (x"ec",x"c2",x"49",x"bf"),
  1874 => (x"a1",x"c1",x"48",x"f0"),
  1875 => (x"b7",x"c0",x"c4",x"78"),
  1876 => (x"87",x"db",x"03",x"a9"),
  1877 => (x"c2",x"48",x"d4",x"ff"),
  1878 => (x"78",x"bf",x"f4",x"ec"),
  1879 => (x"bf",x"f0",x"ec",x"c2"),
  1880 => (x"f0",x"ec",x"c2",x"49"),
  1881 => (x"78",x"a1",x"c1",x"48"),
  1882 => (x"a9",x"b7",x"c0",x"c4"),
  1883 => (x"ff",x"87",x"e5",x"04"),
  1884 => (x"78",x"c8",x"48",x"d0"),
  1885 => (x"48",x"fc",x"ec",x"c2"),
  1886 => (x"4f",x"26",x"78",x"c0"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"5f",x"00",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"5f"),
  1891 => (x"00",x"03",x"03",x"00"),
  1892 => (x"00",x"00",x"03",x"03"),
  1893 => (x"14",x"7f",x"7f",x"14"),
  1894 => (x"00",x"14",x"7f",x"7f"),
  1895 => (x"6b",x"2e",x"24",x"00"),
  1896 => (x"00",x"12",x"3a",x"6b"),
  1897 => (x"18",x"36",x"6a",x"4c"),
  1898 => (x"00",x"32",x"56",x"6c"),
  1899 => (x"59",x"4f",x"7e",x"30"),
  1900 => (x"40",x"68",x"3a",x"77"),
  1901 => (x"07",x"04",x"00",x"00"),
  1902 => (x"00",x"00",x"00",x"03"),
  1903 => (x"3e",x"1c",x"00",x"00"),
  1904 => (x"00",x"00",x"41",x"63"),
  1905 => (x"63",x"41",x"00",x"00"),
  1906 => (x"00",x"00",x"1c",x"3e"),
  1907 => (x"1c",x"3e",x"2a",x"08"),
  1908 => (x"08",x"2a",x"3e",x"1c"),
  1909 => (x"3e",x"08",x"08",x"00"),
  1910 => (x"00",x"08",x"08",x"3e"),
  1911 => (x"e0",x"80",x"00",x"00"),
  1912 => (x"00",x"00",x"00",x"60"),
  1913 => (x"08",x"08",x"08",x"00"),
  1914 => (x"00",x"08",x"08",x"08"),
  1915 => (x"60",x"00",x"00",x"00"),
  1916 => (x"00",x"00",x"00",x"60"),
  1917 => (x"18",x"30",x"60",x"40"),
  1918 => (x"01",x"03",x"06",x"0c"),
  1919 => (x"59",x"7f",x"3e",x"00"),
  1920 => (x"00",x"3e",x"7f",x"4d"),
  1921 => (x"7f",x"06",x"04",x"00"),
  1922 => (x"00",x"00",x"00",x"7f"),
  1923 => (x"71",x"63",x"42",x"00"),
  1924 => (x"00",x"46",x"4f",x"59"),
  1925 => (x"49",x"63",x"22",x"00"),
  1926 => (x"00",x"36",x"7f",x"49"),
  1927 => (x"13",x"16",x"1c",x"18"),
  1928 => (x"00",x"10",x"7f",x"7f"),
  1929 => (x"45",x"67",x"27",x"00"),
  1930 => (x"00",x"39",x"7d",x"45"),
  1931 => (x"4b",x"7e",x"3c",x"00"),
  1932 => (x"00",x"30",x"79",x"49"),
  1933 => (x"71",x"01",x"01",x"00"),
  1934 => (x"00",x"07",x"0f",x"79"),
  1935 => (x"49",x"7f",x"36",x"00"),
  1936 => (x"00",x"36",x"7f",x"49"),
  1937 => (x"49",x"4f",x"06",x"00"),
  1938 => (x"00",x"1e",x"3f",x"69"),
  1939 => (x"66",x"00",x"00",x"00"),
  1940 => (x"00",x"00",x"00",x"66"),
  1941 => (x"e6",x"80",x"00",x"00"),
  1942 => (x"00",x"00",x"00",x"66"),
  1943 => (x"14",x"08",x"08",x"00"),
  1944 => (x"00",x"22",x"22",x"14"),
  1945 => (x"14",x"14",x"14",x"00"),
  1946 => (x"00",x"14",x"14",x"14"),
  1947 => (x"14",x"22",x"22",x"00"),
  1948 => (x"00",x"08",x"08",x"14"),
  1949 => (x"51",x"03",x"02",x"00"),
  1950 => (x"00",x"06",x"0f",x"59"),
  1951 => (x"5d",x"41",x"7f",x"3e"),
  1952 => (x"00",x"1e",x"1f",x"55"),
  1953 => (x"09",x"7f",x"7e",x"00"),
  1954 => (x"00",x"7e",x"7f",x"09"),
  1955 => (x"49",x"7f",x"7f",x"00"),
  1956 => (x"00",x"36",x"7f",x"49"),
  1957 => (x"63",x"3e",x"1c",x"00"),
  1958 => (x"00",x"41",x"41",x"41"),
  1959 => (x"41",x"7f",x"7f",x"00"),
  1960 => (x"00",x"1c",x"3e",x"63"),
  1961 => (x"49",x"7f",x"7f",x"00"),
  1962 => (x"00",x"41",x"41",x"49"),
  1963 => (x"09",x"7f",x"7f",x"00"),
  1964 => (x"00",x"01",x"01",x"09"),
  1965 => (x"41",x"7f",x"3e",x"00"),
  1966 => (x"00",x"7a",x"7b",x"49"),
  1967 => (x"08",x"7f",x"7f",x"00"),
  1968 => (x"00",x"7f",x"7f",x"08"),
  1969 => (x"7f",x"41",x"00",x"00"),
  1970 => (x"00",x"00",x"41",x"7f"),
  1971 => (x"40",x"60",x"20",x"00"),
  1972 => (x"00",x"3f",x"7f",x"40"),
  1973 => (x"1c",x"08",x"7f",x"7f"),
  1974 => (x"00",x"41",x"63",x"36"),
  1975 => (x"40",x"7f",x"7f",x"00"),
  1976 => (x"00",x"40",x"40",x"40"),
  1977 => (x"0c",x"06",x"7f",x"7f"),
  1978 => (x"00",x"7f",x"7f",x"06"),
  1979 => (x"0c",x"06",x"7f",x"7f"),
  1980 => (x"00",x"7f",x"7f",x"18"),
  1981 => (x"41",x"7f",x"3e",x"00"),
  1982 => (x"00",x"3e",x"7f",x"41"),
  1983 => (x"09",x"7f",x"7f",x"00"),
  1984 => (x"00",x"06",x"0f",x"09"),
  1985 => (x"61",x"41",x"7f",x"3e"),
  1986 => (x"00",x"40",x"7e",x"7f"),
  1987 => (x"09",x"7f",x"7f",x"00"),
  1988 => (x"00",x"66",x"7f",x"19"),
  1989 => (x"4d",x"6f",x"26",x"00"),
  1990 => (x"00",x"32",x"7b",x"59"),
  1991 => (x"7f",x"01",x"01",x"00"),
  1992 => (x"00",x"01",x"01",x"7f"),
  1993 => (x"40",x"7f",x"3f",x"00"),
  1994 => (x"00",x"3f",x"7f",x"40"),
  1995 => (x"70",x"3f",x"0f",x"00"),
  1996 => (x"00",x"0f",x"3f",x"70"),
  1997 => (x"18",x"30",x"7f",x"7f"),
  1998 => (x"00",x"7f",x"7f",x"30"),
  1999 => (x"1c",x"36",x"63",x"41"),
  2000 => (x"41",x"63",x"36",x"1c"),
  2001 => (x"7c",x"06",x"03",x"01"),
  2002 => (x"01",x"03",x"06",x"7c"),
  2003 => (x"4d",x"59",x"71",x"61"),
  2004 => (x"00",x"41",x"43",x"47"),
  2005 => (x"7f",x"7f",x"00",x"00"),
  2006 => (x"00",x"00",x"41",x"41"),
  2007 => (x"0c",x"06",x"03",x"01"),
  2008 => (x"40",x"60",x"30",x"18"),
  2009 => (x"41",x"41",x"00",x"00"),
  2010 => (x"00",x"00",x"7f",x"7f"),
  2011 => (x"03",x"06",x"0c",x"08"),
  2012 => (x"00",x"08",x"0c",x"06"),
  2013 => (x"80",x"80",x"80",x"80"),
  2014 => (x"00",x"80",x"80",x"80"),
  2015 => (x"03",x"00",x"00",x"00"),
  2016 => (x"00",x"00",x"04",x"07"),
  2017 => (x"54",x"74",x"20",x"00"),
  2018 => (x"00",x"78",x"7c",x"54"),
  2019 => (x"44",x"7f",x"7f",x"00"),
  2020 => (x"00",x"38",x"7c",x"44"),
  2021 => (x"44",x"7c",x"38",x"00"),
  2022 => (x"00",x"00",x"44",x"44"),
  2023 => (x"44",x"7c",x"38",x"00"),
  2024 => (x"00",x"7f",x"7f",x"44"),
  2025 => (x"54",x"7c",x"38",x"00"),
  2026 => (x"00",x"18",x"5c",x"54"),
  2027 => (x"7f",x"7e",x"04",x"00"),
  2028 => (x"00",x"00",x"05",x"05"),
  2029 => (x"a4",x"bc",x"18",x"00"),
  2030 => (x"00",x"7c",x"fc",x"a4"),
  2031 => (x"04",x"7f",x"7f",x"00"),
  2032 => (x"00",x"78",x"7c",x"04"),
  2033 => (x"3d",x"00",x"00",x"00"),
  2034 => (x"00",x"00",x"40",x"7d"),
  2035 => (x"80",x"80",x"80",x"00"),
  2036 => (x"00",x"00",x"7d",x"fd"),
  2037 => (x"10",x"7f",x"7f",x"00"),
  2038 => (x"00",x"44",x"6c",x"38"),
  2039 => (x"3f",x"00",x"00",x"00"),
  2040 => (x"00",x"00",x"40",x"7f"),
  2041 => (x"18",x"0c",x"7c",x"7c"),
  2042 => (x"00",x"78",x"7c",x"0c"),
  2043 => (x"04",x"7c",x"7c",x"00"),
  2044 => (x"00",x"78",x"7c",x"04"),
  2045 => (x"44",x"7c",x"38",x"00"),
  2046 => (x"00",x"38",x"7c",x"44"),
  2047 => (x"24",x"fc",x"fc",x"00"),
  2048 => (x"00",x"18",x"3c",x"24"),
  2049 => (x"24",x"3c",x"18",x"00"),
  2050 => (x"00",x"fc",x"fc",x"24"),
  2051 => (x"04",x"7c",x"7c",x"00"),
  2052 => (x"00",x"08",x"0c",x"04"),
  2053 => (x"54",x"5c",x"48",x"00"),
  2054 => (x"00",x"20",x"74",x"54"),
  2055 => (x"7f",x"3f",x"04",x"00"),
  2056 => (x"00",x"00",x"44",x"44"),
  2057 => (x"40",x"7c",x"3c",x"00"),
  2058 => (x"00",x"7c",x"7c",x"40"),
  2059 => (x"60",x"3c",x"1c",x"00"),
  2060 => (x"00",x"1c",x"3c",x"60"),
  2061 => (x"30",x"60",x"7c",x"3c"),
  2062 => (x"00",x"3c",x"7c",x"60"),
  2063 => (x"10",x"38",x"6c",x"44"),
  2064 => (x"00",x"44",x"6c",x"38"),
  2065 => (x"e0",x"bc",x"1c",x"00"),
  2066 => (x"00",x"1c",x"3c",x"60"),
  2067 => (x"74",x"64",x"44",x"00"),
  2068 => (x"00",x"44",x"4c",x"5c"),
  2069 => (x"3e",x"08",x"08",x"00"),
  2070 => (x"00",x"41",x"41",x"77"),
  2071 => (x"7f",x"00",x"00",x"00"),
  2072 => (x"00",x"00",x"00",x"7f"),
  2073 => (x"77",x"41",x"41",x"00"),
  2074 => (x"00",x"08",x"08",x"3e"),
  2075 => (x"03",x"01",x"01",x"02"),
  2076 => (x"00",x"01",x"02",x"02"),
  2077 => (x"7f",x"7f",x"7f",x"7f"),
  2078 => (x"00",x"7f",x"7f",x"7f"),
  2079 => (x"1c",x"1c",x"08",x"08"),
  2080 => (x"7f",x"7f",x"3e",x"3e"),
  2081 => (x"3e",x"3e",x"7f",x"7f"),
  2082 => (x"08",x"08",x"1c",x"1c"),
  2083 => (x"7c",x"18",x"10",x"00"),
  2084 => (x"00",x"10",x"18",x"7c"),
  2085 => (x"7c",x"30",x"10",x"00"),
  2086 => (x"00",x"10",x"30",x"7c"),
  2087 => (x"60",x"60",x"30",x"10"),
  2088 => (x"00",x"06",x"1e",x"78"),
  2089 => (x"18",x"3c",x"66",x"42"),
  2090 => (x"00",x"42",x"66",x"3c"),
  2091 => (x"c2",x"6a",x"38",x"78"),
  2092 => (x"00",x"38",x"6c",x"c6"),
  2093 => (x"60",x"00",x"00",x"60"),
  2094 => (x"00",x"60",x"00",x"00"),
  2095 => (x"5c",x"5b",x"5e",x"0e"),
  2096 => (x"71",x"1e",x"0e",x"5d"),
  2097 => (x"c1",x"ed",x"c2",x"4c"),
  2098 => (x"4b",x"c0",x"4d",x"bf"),
  2099 => (x"ab",x"74",x"1e",x"c0"),
  2100 => (x"c4",x"87",x"c7",x"02"),
  2101 => (x"78",x"c0",x"48",x"a6"),
  2102 => (x"a6",x"c4",x"87",x"c5"),
  2103 => (x"c4",x"78",x"c1",x"48"),
  2104 => (x"49",x"73",x"1e",x"66"),
  2105 => (x"c8",x"87",x"df",x"ee"),
  2106 => (x"49",x"e0",x"c0",x"86"),
  2107 => (x"c4",x"87",x"ee",x"ef"),
  2108 => (x"49",x"6a",x"4a",x"a5"),
  2109 => (x"f1",x"87",x"f0",x"f0"),
  2110 => (x"85",x"cb",x"87",x"c6"),
  2111 => (x"b7",x"c8",x"83",x"c1"),
  2112 => (x"c7",x"ff",x"04",x"ab"),
  2113 => (x"4d",x"26",x"26",x"87"),
  2114 => (x"4b",x"26",x"4c",x"26"),
  2115 => (x"71",x"1e",x"4f",x"26"),
  2116 => (x"c5",x"ed",x"c2",x"4a"),
  2117 => (x"c5",x"ed",x"c2",x"5a"),
  2118 => (x"49",x"78",x"c7",x"48"),
  2119 => (x"26",x"87",x"dd",x"fe"),
  2120 => (x"1e",x"73",x"1e",x"4f"),
  2121 => (x"b7",x"c0",x"4a",x"71"),
  2122 => (x"87",x"d3",x"03",x"aa"),
  2123 => (x"bf",x"db",x"d3",x"c2"),
  2124 => (x"c1",x"87",x"c4",x"05"),
  2125 => (x"c0",x"87",x"c2",x"4b"),
  2126 => (x"df",x"d3",x"c2",x"4b"),
  2127 => (x"c2",x"87",x"c4",x"5b"),
  2128 => (x"c2",x"5a",x"df",x"d3"),
  2129 => (x"4a",x"bf",x"db",x"d3"),
  2130 => (x"c0",x"c1",x"9a",x"c1"),
  2131 => (x"e8",x"ec",x"49",x"a2"),
  2132 => (x"c2",x"48",x"fc",x"87"),
  2133 => (x"78",x"bf",x"db",x"d3"),
  2134 => (x"1e",x"87",x"ef",x"fe"),
  2135 => (x"66",x"c4",x"4a",x"71"),
  2136 => (x"ea",x"49",x"72",x"1e"),
  2137 => (x"26",x"26",x"87",x"ee"),
  2138 => (x"d4",x"ff",x"1e",x"4f"),
  2139 => (x"78",x"ff",x"c3",x"48"),
  2140 => (x"c0",x"48",x"d0",x"ff"),
  2141 => (x"d4",x"ff",x"78",x"e1"),
  2142 => (x"71",x"78",x"c1",x"48"),
  2143 => (x"ff",x"30",x"c4",x"48"),
  2144 => (x"ff",x"78",x"08",x"d4"),
  2145 => (x"e0",x"c0",x"48",x"d0"),
  2146 => (x"0e",x"4f",x"26",x"78"),
  2147 => (x"5d",x"5c",x"5b",x"5e"),
  2148 => (x"c4",x"86",x"f4",x"0e"),
  2149 => (x"78",x"c0",x"48",x"a6"),
  2150 => (x"7e",x"bf",x"ec",x"4b"),
  2151 => (x"bf",x"c1",x"ed",x"c2"),
  2152 => (x"4c",x"bf",x"e8",x"4d"),
  2153 => (x"bf",x"db",x"d3",x"c2"),
  2154 => (x"87",x"d6",x"e2",x"49"),
  2155 => (x"cc",x"49",x"ee",x"cb"),
  2156 => (x"a6",x"cc",x"87",x"f1"),
  2157 => (x"e6",x"49",x"c7",x"58"),
  2158 => (x"98",x"70",x"87",x"cb"),
  2159 => (x"6e",x"87",x"c8",x"05"),
  2160 => (x"02",x"99",x"c1",x"49"),
  2161 => (x"c1",x"87",x"c3",x"c1"),
  2162 => (x"7e",x"bf",x"ec",x"4b"),
  2163 => (x"bf",x"db",x"d3",x"c2"),
  2164 => (x"87",x"ee",x"e1",x"49"),
  2165 => (x"cc",x"49",x"66",x"c8"),
  2166 => (x"98",x"70",x"87",x"d5"),
  2167 => (x"c2",x"87",x"d8",x"02"),
  2168 => (x"49",x"bf",x"d3",x"d3"),
  2169 => (x"d3",x"c2",x"b9",x"c1"),
  2170 => (x"fd",x"71",x"59",x"d7"),
  2171 => (x"ee",x"cb",x"87",x"fb"),
  2172 => (x"87",x"ef",x"cb",x"49"),
  2173 => (x"c7",x"58",x"a6",x"cc"),
  2174 => (x"87",x"c9",x"e5",x"49"),
  2175 => (x"ff",x"05",x"98",x"70"),
  2176 => (x"49",x"6e",x"87",x"c5"),
  2177 => (x"fe",x"05",x"99",x"c1"),
  2178 => (x"9b",x"73",x"87",x"fd"),
  2179 => (x"ff",x"87",x"d0",x"02"),
  2180 => (x"87",x"cd",x"fc",x"49"),
  2181 => (x"e4",x"49",x"da",x"c1"),
  2182 => (x"a6",x"c4",x"87",x"eb"),
  2183 => (x"c2",x"78",x"c1",x"48"),
  2184 => (x"05",x"bf",x"db",x"d3"),
  2185 => (x"c3",x"87",x"e9",x"c0"),
  2186 => (x"d8",x"e4",x"49",x"fd"),
  2187 => (x"49",x"fa",x"c3",x"87"),
  2188 => (x"74",x"87",x"d2",x"e4"),
  2189 => (x"99",x"ff",x"c3",x"49"),
  2190 => (x"49",x"c0",x"1e",x"71"),
  2191 => (x"74",x"87",x"dc",x"fc"),
  2192 => (x"29",x"b7",x"c8",x"49"),
  2193 => (x"49",x"c1",x"1e",x"71"),
  2194 => (x"c8",x"87",x"d0",x"fc"),
  2195 => (x"87",x"ed",x"c8",x"86"),
  2196 => (x"ff",x"c3",x"49",x"74"),
  2197 => (x"2c",x"b7",x"c8",x"99"),
  2198 => (x"9c",x"74",x"b4",x"71"),
  2199 => (x"c2",x"87",x"dd",x"02"),
  2200 => (x"49",x"bf",x"d7",x"d3"),
  2201 => (x"70",x"87",x"c8",x"ca"),
  2202 => (x"87",x"c4",x"05",x"98"),
  2203 => (x"87",x"d2",x"4c",x"c0"),
  2204 => (x"c9",x"49",x"e0",x"c2"),
  2205 => (x"d3",x"c2",x"87",x"ed"),
  2206 => (x"87",x"c6",x"58",x"db"),
  2207 => (x"48",x"d7",x"d3",x"c2"),
  2208 => (x"49",x"74",x"78",x"c0"),
  2209 => (x"cd",x"05",x"99",x"c2"),
  2210 => (x"49",x"eb",x"c3",x"87"),
  2211 => (x"70",x"87",x"f6",x"e2"),
  2212 => (x"02",x"99",x"c2",x"49"),
  2213 => (x"d8",x"c1",x"87",x"cf"),
  2214 => (x"bf",x"6e",x"7e",x"a5"),
  2215 => (x"87",x"c5",x"c0",x"02"),
  2216 => (x"73",x"49",x"fb",x"4b"),
  2217 => (x"c1",x"49",x"74",x"0f"),
  2218 => (x"87",x"cd",x"05",x"99"),
  2219 => (x"e2",x"49",x"f4",x"c3"),
  2220 => (x"49",x"70",x"87",x"d3"),
  2221 => (x"cf",x"02",x"99",x"c2"),
  2222 => (x"a5",x"d8",x"c1",x"87"),
  2223 => (x"02",x"bf",x"6e",x"7e"),
  2224 => (x"4b",x"87",x"c5",x"c0"),
  2225 => (x"0f",x"73",x"49",x"fa"),
  2226 => (x"99",x"c8",x"49",x"74"),
  2227 => (x"c3",x"87",x"ce",x"05"),
  2228 => (x"f0",x"e1",x"49",x"f5"),
  2229 => (x"c2",x"49",x"70",x"87"),
  2230 => (x"e5",x"c0",x"02",x"99"),
  2231 => (x"c5",x"ed",x"c2",x"87"),
  2232 => (x"ca",x"c0",x"02",x"bf"),
  2233 => (x"88",x"c1",x"48",x"87"),
  2234 => (x"58",x"c9",x"ed",x"c2"),
  2235 => (x"c1",x"87",x"ce",x"c0"),
  2236 => (x"6a",x"4a",x"a5",x"d8"),
  2237 => (x"87",x"c5",x"c0",x"02"),
  2238 => (x"73",x"49",x"ff",x"4b"),
  2239 => (x"48",x"a6",x"c4",x"0f"),
  2240 => (x"49",x"74",x"78",x"c1"),
  2241 => (x"c0",x"05",x"99",x"c4"),
  2242 => (x"f2",x"c3",x"87",x"ce"),
  2243 => (x"87",x"f5",x"e0",x"49"),
  2244 => (x"99",x"c2",x"49",x"70"),
  2245 => (x"87",x"ec",x"c0",x"02"),
  2246 => (x"bf",x"c5",x"ed",x"c2"),
  2247 => (x"b7",x"c7",x"48",x"7e"),
  2248 => (x"cb",x"c0",x"03",x"a8"),
  2249 => (x"c1",x"48",x"6e",x"87"),
  2250 => (x"c9",x"ed",x"c2",x"80"),
  2251 => (x"87",x"cf",x"c0",x"58"),
  2252 => (x"7e",x"a5",x"d8",x"c1"),
  2253 => (x"c0",x"02",x"bf",x"6e"),
  2254 => (x"fe",x"4b",x"87",x"c5"),
  2255 => (x"c4",x"0f",x"73",x"49"),
  2256 => (x"78",x"c1",x"48",x"a6"),
  2257 => (x"ff",x"49",x"fd",x"c3"),
  2258 => (x"70",x"87",x"fa",x"df"),
  2259 => (x"02",x"99",x"c2",x"49"),
  2260 => (x"c2",x"87",x"e5",x"c0"),
  2261 => (x"02",x"bf",x"c5",x"ed"),
  2262 => (x"c2",x"87",x"c9",x"c0"),
  2263 => (x"c0",x"48",x"c5",x"ed"),
  2264 => (x"87",x"cf",x"c0",x"78"),
  2265 => (x"7e",x"a5",x"d8",x"c1"),
  2266 => (x"c0",x"02",x"bf",x"6e"),
  2267 => (x"fd",x"4b",x"87",x"c5"),
  2268 => (x"c4",x"0f",x"73",x"49"),
  2269 => (x"78",x"c1",x"48",x"a6"),
  2270 => (x"ff",x"49",x"fa",x"c3"),
  2271 => (x"70",x"87",x"c6",x"df"),
  2272 => (x"02",x"99",x"c2",x"49"),
  2273 => (x"c2",x"87",x"e9",x"c0"),
  2274 => (x"48",x"bf",x"c5",x"ed"),
  2275 => (x"03",x"a8",x"b7",x"c7"),
  2276 => (x"c2",x"87",x"c9",x"c0"),
  2277 => (x"c7",x"48",x"c5",x"ed"),
  2278 => (x"87",x"cf",x"c0",x"78"),
  2279 => (x"7e",x"a5",x"d8",x"c1"),
  2280 => (x"c0",x"02",x"bf",x"6e"),
  2281 => (x"fc",x"4b",x"87",x"c5"),
  2282 => (x"c4",x"0f",x"73",x"49"),
  2283 => (x"78",x"c1",x"48",x"a6"),
  2284 => (x"ed",x"c2",x"4b",x"c0"),
  2285 => (x"50",x"c0",x"48",x"c0"),
  2286 => (x"c4",x"49",x"ee",x"cb"),
  2287 => (x"a6",x"cc",x"87",x"e5"),
  2288 => (x"c0",x"ed",x"c2",x"58"),
  2289 => (x"c1",x"05",x"bf",x"97"),
  2290 => (x"49",x"74",x"87",x"de"),
  2291 => (x"05",x"99",x"f0",x"c3"),
  2292 => (x"c1",x"87",x"cd",x"c0"),
  2293 => (x"dd",x"ff",x"49",x"da"),
  2294 => (x"98",x"70",x"87",x"eb"),
  2295 => (x"87",x"c8",x"c1",x"02"),
  2296 => (x"bf",x"e8",x"4b",x"c1"),
  2297 => (x"ff",x"c3",x"49",x"4c"),
  2298 => (x"2c",x"b7",x"c8",x"99"),
  2299 => (x"d3",x"c2",x"b4",x"71"),
  2300 => (x"ff",x"49",x"bf",x"db"),
  2301 => (x"c8",x"87",x"cb",x"d9"),
  2302 => (x"f2",x"c3",x"49",x"66"),
  2303 => (x"02",x"98",x"70",x"87"),
  2304 => (x"c2",x"87",x"c6",x"c0"),
  2305 => (x"c1",x"48",x"c0",x"ed"),
  2306 => (x"c0",x"ed",x"c2",x"50"),
  2307 => (x"c0",x"05",x"bf",x"97"),
  2308 => (x"49",x"74",x"87",x"d6"),
  2309 => (x"05",x"99",x"f0",x"c3"),
  2310 => (x"c1",x"87",x"c5",x"ff"),
  2311 => (x"dc",x"ff",x"49",x"da"),
  2312 => (x"98",x"70",x"87",x"e3"),
  2313 => (x"87",x"f8",x"fe",x"05"),
  2314 => (x"c0",x"02",x"9b",x"73"),
  2315 => (x"a6",x"c8",x"87",x"dc"),
  2316 => (x"c5",x"ed",x"c2",x"48"),
  2317 => (x"66",x"c8",x"78",x"bf"),
  2318 => (x"75",x"91",x"cb",x"49"),
  2319 => (x"bf",x"6e",x"7e",x"a1"),
  2320 => (x"87",x"c6",x"c0",x"02"),
  2321 => (x"49",x"66",x"c8",x"4b"),
  2322 => (x"66",x"c4",x"0f",x"73"),
  2323 => (x"87",x"c8",x"c0",x"02"),
  2324 => (x"bf",x"c5",x"ed",x"c2"),
  2325 => (x"87",x"e4",x"f1",x"49"),
  2326 => (x"bf",x"df",x"d3",x"c2"),
  2327 => (x"87",x"dd",x"c0",x"02"),
  2328 => (x"87",x"cb",x"c2",x"49"),
  2329 => (x"c0",x"02",x"98",x"70"),
  2330 => (x"ed",x"c2",x"87",x"d3"),
  2331 => (x"f1",x"49",x"bf",x"c5"),
  2332 => (x"49",x"c0",x"87",x"ca"),
  2333 => (x"c2",x"87",x"ea",x"f2"),
  2334 => (x"c0",x"48",x"df",x"d3"),
  2335 => (x"f2",x"8e",x"f4",x"78"),
  2336 => (x"5e",x"0e",x"87",x"c4"),
  2337 => (x"0e",x"5d",x"5c",x"5b"),
  2338 => (x"c2",x"4c",x"71",x"1e"),
  2339 => (x"49",x"bf",x"c1",x"ed"),
  2340 => (x"4d",x"a1",x"cd",x"c1"),
  2341 => (x"69",x"81",x"d1",x"c1"),
  2342 => (x"02",x"9c",x"74",x"7e"),
  2343 => (x"a5",x"c4",x"87",x"cf"),
  2344 => (x"c2",x"7b",x"74",x"4b"),
  2345 => (x"49",x"bf",x"c1",x"ed"),
  2346 => (x"6e",x"87",x"e3",x"f1"),
  2347 => (x"05",x"9c",x"74",x"7b"),
  2348 => (x"4b",x"c0",x"87",x"c4"),
  2349 => (x"4b",x"c1",x"87",x"c2"),
  2350 => (x"e4",x"f1",x"49",x"73"),
  2351 => (x"02",x"66",x"d4",x"87"),
  2352 => (x"de",x"49",x"87",x"c7"),
  2353 => (x"c2",x"4a",x"70",x"87"),
  2354 => (x"c2",x"4a",x"c0",x"87"),
  2355 => (x"26",x"5a",x"e3",x"d3"),
  2356 => (x"00",x"87",x"f3",x"f0"),
  2357 => (x"00",x"00",x"00",x"00"),
  2358 => (x"00",x"00",x"00",x"00"),
  2359 => (x"00",x"00",x"00",x"00"),
  2360 => (x"1e",x"00",x"00",x"00"),
  2361 => (x"c8",x"ff",x"4a",x"71"),
  2362 => (x"a1",x"72",x"49",x"bf"),
  2363 => (x"1e",x"4f",x"26",x"48"),
  2364 => (x"89",x"bf",x"c8",x"ff"),
  2365 => (x"c0",x"c0",x"c0",x"fe"),
  2366 => (x"01",x"a9",x"c0",x"c0"),
  2367 => (x"4a",x"c0",x"87",x"c4"),
  2368 => (x"4a",x"c1",x"87",x"c2"),
  2369 => (x"4f",x"26",x"48",x"72"),
  2370 => (x"5c",x"5b",x"5e",x"0e"),
  2371 => (x"4b",x"71",x"0e",x"5d"),
  2372 => (x"d0",x"4c",x"d4",x"ff"),
  2373 => (x"78",x"c0",x"48",x"66"),
  2374 => (x"da",x"ff",x"49",x"d6"),
  2375 => (x"ff",x"c3",x"87",x"df"),
  2376 => (x"c3",x"49",x"6c",x"7c"),
  2377 => (x"4d",x"71",x"99",x"ff"),
  2378 => (x"99",x"f0",x"c3",x"49"),
  2379 => (x"05",x"a9",x"e0",x"c1"),
  2380 => (x"ff",x"c3",x"87",x"cb"),
  2381 => (x"c3",x"48",x"6c",x"7c"),
  2382 => (x"08",x"66",x"d0",x"98"),
  2383 => (x"7c",x"ff",x"c3",x"78"),
  2384 => (x"c8",x"49",x"4a",x"6c"),
  2385 => (x"7c",x"ff",x"c3",x"31"),
  2386 => (x"b2",x"71",x"4a",x"6c"),
  2387 => (x"31",x"c8",x"49",x"72"),
  2388 => (x"6c",x"7c",x"ff",x"c3"),
  2389 => (x"72",x"b2",x"71",x"4a"),
  2390 => (x"c3",x"31",x"c8",x"49"),
  2391 => (x"4a",x"6c",x"7c",x"ff"),
  2392 => (x"d0",x"ff",x"b2",x"71"),
  2393 => (x"78",x"e0",x"c0",x"48"),
  2394 => (x"c2",x"02",x"9b",x"73"),
  2395 => (x"75",x"7b",x"72",x"87"),
  2396 => (x"26",x"4d",x"26",x"48"),
  2397 => (x"26",x"4b",x"26",x"4c"),
  2398 => (x"4f",x"26",x"1e",x"4f"),
  2399 => (x"5c",x"5b",x"5e",x"0e"),
  2400 => (x"76",x"86",x"f8",x"0e"),
  2401 => (x"49",x"a6",x"c8",x"1e"),
  2402 => (x"c4",x"87",x"fd",x"fd"),
  2403 => (x"6e",x"4b",x"70",x"86"),
  2404 => (x"01",x"a8",x"c0",x"48"),
  2405 => (x"73",x"87",x"f0",x"c2"),
  2406 => (x"9a",x"f0",x"c3",x"4a"),
  2407 => (x"02",x"aa",x"d0",x"c1"),
  2408 => (x"e0",x"c1",x"87",x"c7"),
  2409 => (x"de",x"c2",x"05",x"aa"),
  2410 => (x"c8",x"49",x"73",x"87"),
  2411 => (x"87",x"c3",x"02",x"99"),
  2412 => (x"73",x"87",x"c6",x"ff"),
  2413 => (x"c2",x"9c",x"c3",x"4c"),
  2414 => (x"c2",x"c1",x"05",x"ac"),
  2415 => (x"49",x"66",x"c4",x"87"),
  2416 => (x"1e",x"71",x"31",x"c9"),
  2417 => (x"d4",x"4a",x"66",x"c4"),
  2418 => (x"c9",x"ed",x"c2",x"92"),
  2419 => (x"fe",x"81",x"72",x"49"),
  2420 => (x"d8",x"87",x"f4",x"cf"),
  2421 => (x"e4",x"d7",x"ff",x"49"),
  2422 => (x"1e",x"c0",x"c8",x"87"),
  2423 => (x"49",x"f2",x"db",x"c2"),
  2424 => (x"87",x"fa",x"eb",x"fd"),
  2425 => (x"c0",x"48",x"d0",x"ff"),
  2426 => (x"db",x"c2",x"78",x"e0"),
  2427 => (x"66",x"cc",x"1e",x"f2"),
  2428 => (x"c2",x"92",x"d4",x"4a"),
  2429 => (x"72",x"49",x"c9",x"ed"),
  2430 => (x"fc",x"cd",x"fe",x"81"),
  2431 => (x"c1",x"86",x"cc",x"87"),
  2432 => (x"c2",x"c1",x"05",x"ac"),
  2433 => (x"49",x"66",x"c4",x"87"),
  2434 => (x"1e",x"71",x"31",x"c9"),
  2435 => (x"d4",x"4a",x"66",x"c4"),
  2436 => (x"c9",x"ed",x"c2",x"92"),
  2437 => (x"fe",x"81",x"72",x"49"),
  2438 => (x"c2",x"87",x"ec",x"ce"),
  2439 => (x"c8",x"1e",x"f2",x"db"),
  2440 => (x"92",x"d4",x"4a",x"66"),
  2441 => (x"49",x"c9",x"ed",x"c2"),
  2442 => (x"cb",x"fe",x"81",x"72"),
  2443 => (x"49",x"d7",x"87",x"fd"),
  2444 => (x"87",x"c9",x"d6",x"ff"),
  2445 => (x"c2",x"1e",x"c0",x"c8"),
  2446 => (x"fd",x"49",x"f2",x"db"),
  2447 => (x"cc",x"87",x"f8",x"e9"),
  2448 => (x"48",x"d0",x"ff",x"86"),
  2449 => (x"f8",x"78",x"e0",x"c0"),
  2450 => (x"87",x"e7",x"fc",x"8e"),
  2451 => (x"5c",x"5b",x"5e",x"0e"),
  2452 => (x"4a",x"71",x"0e",x"5d"),
  2453 => (x"d0",x"4c",x"d4",x"ff"),
  2454 => (x"b7",x"c3",x"4d",x"66"),
  2455 => (x"87",x"c5",x"06",x"ad"),
  2456 => (x"e1",x"c1",x"48",x"c0"),
  2457 => (x"75",x"1e",x"72",x"87"),
  2458 => (x"c2",x"93",x"d4",x"4b"),
  2459 => (x"73",x"83",x"c9",x"ed"),
  2460 => (x"c4",x"c6",x"fe",x"49"),
  2461 => (x"6b",x"83",x"c8",x"87"),
  2462 => (x"48",x"d0",x"ff",x"4b"),
  2463 => (x"dd",x"78",x"e1",x"c8"),
  2464 => (x"c3",x"48",x"73",x"7c"),
  2465 => (x"7c",x"70",x"98",x"ff"),
  2466 => (x"b7",x"c8",x"49",x"73"),
  2467 => (x"c3",x"48",x"71",x"29"),
  2468 => (x"7c",x"70",x"98",x"ff"),
  2469 => (x"b7",x"d0",x"49",x"73"),
  2470 => (x"c3",x"48",x"71",x"29"),
  2471 => (x"7c",x"70",x"98",x"ff"),
  2472 => (x"b7",x"d8",x"48",x"73"),
  2473 => (x"c0",x"7c",x"70",x"28"),
  2474 => (x"7c",x"7c",x"7c",x"7c"),
  2475 => (x"7c",x"7c",x"7c",x"7c"),
  2476 => (x"7c",x"7c",x"7c",x"7c"),
  2477 => (x"c0",x"48",x"d0",x"ff"),
  2478 => (x"1e",x"75",x"78",x"e0"),
  2479 => (x"d4",x"ff",x"49",x"dc"),
  2480 => (x"86",x"c8",x"87",x"e0"),
  2481 => (x"e8",x"fa",x"48",x"73"),
  2482 => (x"e8",x"fa",x"48",x"87"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

