
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"18",x"3c",x"24"),
     1 => (x"24",x"3c",x"18",x"00"),
     2 => (x"00",x"fc",x"fc",x"24"),
     3 => (x"04",x"7c",x"7c",x"00"),
     4 => (x"00",x"08",x"0c",x"04"),
     5 => (x"54",x"5c",x"48",x"00"),
     6 => (x"00",x"20",x"74",x"54"),
     7 => (x"7f",x"3f",x"04",x"00"),
     8 => (x"00",x"00",x"44",x"44"),
     9 => (x"40",x"7c",x"3c",x"00"),
    10 => (x"00",x"7c",x"7c",x"40"),
    11 => (x"60",x"3c",x"1c",x"00"),
    12 => (x"00",x"1c",x"3c",x"60"),
    13 => (x"30",x"60",x"7c",x"3c"),
    14 => (x"00",x"3c",x"7c",x"60"),
    15 => (x"10",x"38",x"6c",x"44"),
    16 => (x"00",x"44",x"6c",x"38"),
    17 => (x"e0",x"bc",x"1c",x"00"),
    18 => (x"00",x"1c",x"3c",x"60"),
    19 => (x"74",x"64",x"44",x"00"),
    20 => (x"00",x"44",x"4c",x"5c"),
    21 => (x"3e",x"08",x"08",x"00"),
    22 => (x"00",x"41",x"41",x"77"),
    23 => (x"7f",x"00",x"00",x"00"),
    24 => (x"00",x"00",x"00",x"7f"),
    25 => (x"77",x"41",x"41",x"00"),
    26 => (x"00",x"08",x"08",x"3e"),
    27 => (x"03",x"01",x"01",x"02"),
    28 => (x"00",x"01",x"02",x"02"),
    29 => (x"7f",x"7f",x"7f",x"7f"),
    30 => (x"00",x"7f",x"7f",x"7f"),
    31 => (x"1c",x"1c",x"08",x"08"),
    32 => (x"7f",x"7f",x"3e",x"3e"),
    33 => (x"3e",x"3e",x"7f",x"7f"),
    34 => (x"08",x"08",x"1c",x"1c"),
    35 => (x"7c",x"18",x"10",x"00"),
    36 => (x"00",x"10",x"18",x"7c"),
    37 => (x"7c",x"30",x"10",x"00"),
    38 => (x"00",x"10",x"30",x"7c"),
    39 => (x"60",x"60",x"30",x"10"),
    40 => (x"00",x"06",x"1e",x"78"),
    41 => (x"18",x"3c",x"66",x"42"),
    42 => (x"00",x"42",x"66",x"3c"),
    43 => (x"c2",x"6a",x"38",x"78"),
    44 => (x"00",x"38",x"6c",x"c6"),
    45 => (x"60",x"00",x"00",x"60"),
    46 => (x"00",x"60",x"00",x"00"),
    47 => (x"5c",x"5b",x"5e",x"0e"),
    48 => (x"71",x"1e",x"0e",x"5d"),
    49 => (x"c1",x"ed",x"c2",x"4c"),
    50 => (x"4b",x"c0",x"4d",x"bf"),
    51 => (x"ab",x"74",x"1e",x"c0"),
    52 => (x"c4",x"87",x"c7",x"02"),
    53 => (x"78",x"c0",x"48",x"a6"),
    54 => (x"a6",x"c4",x"87",x"c5"),
    55 => (x"c4",x"78",x"c1",x"48"),
    56 => (x"49",x"73",x"1e",x"66"),
    57 => (x"c8",x"87",x"df",x"ee"),
    58 => (x"49",x"e0",x"c0",x"86"),
    59 => (x"c4",x"87",x"ee",x"ef"),
    60 => (x"49",x"6a",x"4a",x"a5"),
    61 => (x"f1",x"87",x"f0",x"f0"),
    62 => (x"85",x"cb",x"87",x"c6"),
    63 => (x"b7",x"c8",x"83",x"c1"),
    64 => (x"c7",x"ff",x"04",x"ab"),
    65 => (x"4d",x"26",x"26",x"87"),
    66 => (x"4b",x"26",x"4c",x"26"),
    67 => (x"71",x"1e",x"4f",x"26"),
    68 => (x"c5",x"ed",x"c2",x"4a"),
    69 => (x"c5",x"ed",x"c2",x"5a"),
    70 => (x"49",x"78",x"c7",x"48"),
    71 => (x"26",x"87",x"dd",x"fe"),
    72 => (x"1e",x"73",x"1e",x"4f"),
    73 => (x"b7",x"c0",x"4a",x"71"),
    74 => (x"87",x"d3",x"03",x"aa"),
    75 => (x"bf",x"db",x"d3",x"c2"),
    76 => (x"c1",x"87",x"c4",x"05"),
    77 => (x"c0",x"87",x"c2",x"4b"),
    78 => (x"df",x"d3",x"c2",x"4b"),
    79 => (x"c2",x"87",x"c4",x"5b"),
    80 => (x"c2",x"5a",x"df",x"d3"),
    81 => (x"4a",x"bf",x"db",x"d3"),
    82 => (x"c0",x"c1",x"9a",x"c1"),
    83 => (x"e8",x"ec",x"49",x"a2"),
    84 => (x"c2",x"48",x"fc",x"87"),
    85 => (x"78",x"bf",x"db",x"d3"),
    86 => (x"1e",x"87",x"ef",x"fe"),
    87 => (x"66",x"c4",x"4a",x"71"),
    88 => (x"ea",x"49",x"72",x"1e"),
    89 => (x"26",x"26",x"87",x"ee"),
    90 => (x"d4",x"ff",x"1e",x"4f"),
    91 => (x"78",x"ff",x"c3",x"48"),
    92 => (x"c0",x"48",x"d0",x"ff"),
    93 => (x"d4",x"ff",x"78",x"e1"),
    94 => (x"71",x"78",x"c1",x"48"),
    95 => (x"ff",x"30",x"c4",x"48"),
    96 => (x"ff",x"78",x"08",x"d4"),
    97 => (x"e0",x"c0",x"48",x"d0"),
    98 => (x"0e",x"4f",x"26",x"78"),
    99 => (x"5d",x"5c",x"5b",x"5e"),
   100 => (x"c4",x"86",x"f4",x"0e"),
   101 => (x"78",x"c0",x"48",x"a6"),
   102 => (x"7e",x"bf",x"ec",x"4b"),
   103 => (x"bf",x"c1",x"ed",x"c2"),
   104 => (x"4c",x"bf",x"e8",x"4d"),
   105 => (x"bf",x"db",x"d3",x"c2"),
   106 => (x"87",x"d6",x"e2",x"49"),
   107 => (x"cc",x"49",x"ee",x"cb"),
   108 => (x"a6",x"cc",x"87",x"f1"),
   109 => (x"e6",x"49",x"c7",x"58"),
   110 => (x"98",x"70",x"87",x"cb"),
   111 => (x"6e",x"87",x"c8",x"05"),
   112 => (x"02",x"99",x"c1",x"49"),
   113 => (x"c1",x"87",x"c3",x"c1"),
   114 => (x"7e",x"bf",x"ec",x"4b"),
   115 => (x"bf",x"db",x"d3",x"c2"),
   116 => (x"87",x"ee",x"e1",x"49"),
   117 => (x"cc",x"49",x"66",x"c8"),
   118 => (x"98",x"70",x"87",x"d5"),
   119 => (x"c2",x"87",x"d8",x"02"),
   120 => (x"49",x"bf",x"d3",x"d3"),
   121 => (x"d3",x"c2",x"b9",x"c1"),
   122 => (x"fd",x"71",x"59",x"d7"),
   123 => (x"ee",x"cb",x"87",x"fb"),
   124 => (x"87",x"ef",x"cb",x"49"),
   125 => (x"c7",x"58",x"a6",x"cc"),
   126 => (x"87",x"c9",x"e5",x"49"),
   127 => (x"ff",x"05",x"98",x"70"),
   128 => (x"49",x"6e",x"87",x"c5"),
   129 => (x"fe",x"05",x"99",x"c1"),
   130 => (x"9b",x"73",x"87",x"fd"),
   131 => (x"ff",x"87",x"d0",x"02"),
   132 => (x"87",x"cd",x"fc",x"49"),
   133 => (x"e4",x"49",x"da",x"c1"),
   134 => (x"a6",x"c4",x"87",x"eb"),
   135 => (x"c2",x"78",x"c1",x"48"),
   136 => (x"05",x"bf",x"db",x"d3"),
   137 => (x"c3",x"87",x"e9",x"c0"),
   138 => (x"d8",x"e4",x"49",x"fd"),
   139 => (x"49",x"fa",x"c3",x"87"),
   140 => (x"74",x"87",x"d2",x"e4"),
   141 => (x"99",x"ff",x"c3",x"49"),
   142 => (x"49",x"c0",x"1e",x"71"),
   143 => (x"74",x"87",x"dc",x"fc"),
   144 => (x"29",x"b7",x"c8",x"49"),
   145 => (x"49",x"c1",x"1e",x"71"),
   146 => (x"c8",x"87",x"d0",x"fc"),
   147 => (x"87",x"ed",x"c8",x"86"),
   148 => (x"ff",x"c3",x"49",x"74"),
   149 => (x"2c",x"b7",x"c8",x"99"),
   150 => (x"9c",x"74",x"b4",x"71"),
   151 => (x"c2",x"87",x"dd",x"02"),
   152 => (x"49",x"bf",x"d7",x"d3"),
   153 => (x"70",x"87",x"c8",x"ca"),
   154 => (x"87",x"c4",x"05",x"98"),
   155 => (x"87",x"d2",x"4c",x"c0"),
   156 => (x"c9",x"49",x"e0",x"c2"),
   157 => (x"d3",x"c2",x"87",x"ed"),
   158 => (x"87",x"c6",x"58",x"db"),
   159 => (x"48",x"d7",x"d3",x"c2"),
   160 => (x"49",x"74",x"78",x"c0"),
   161 => (x"cd",x"05",x"99",x"c2"),
   162 => (x"49",x"eb",x"c3",x"87"),
   163 => (x"70",x"87",x"f6",x"e2"),
   164 => (x"02",x"99",x"c2",x"49"),
   165 => (x"d8",x"c1",x"87",x"cf"),
   166 => (x"bf",x"6e",x"7e",x"a5"),
   167 => (x"87",x"c5",x"c0",x"02"),
   168 => (x"73",x"49",x"fb",x"4b"),
   169 => (x"c1",x"49",x"74",x"0f"),
   170 => (x"87",x"cd",x"05",x"99"),
   171 => (x"e2",x"49",x"f4",x"c3"),
   172 => (x"49",x"70",x"87",x"d3"),
   173 => (x"cf",x"02",x"99",x"c2"),
   174 => (x"a5",x"d8",x"c1",x"87"),
   175 => (x"02",x"bf",x"6e",x"7e"),
   176 => (x"4b",x"87",x"c5",x"c0"),
   177 => (x"0f",x"73",x"49",x"fa"),
   178 => (x"99",x"c8",x"49",x"74"),
   179 => (x"c3",x"87",x"ce",x"05"),
   180 => (x"f0",x"e1",x"49",x"f5"),
   181 => (x"c2",x"49",x"70",x"87"),
   182 => (x"e5",x"c0",x"02",x"99"),
   183 => (x"c5",x"ed",x"c2",x"87"),
   184 => (x"ca",x"c0",x"02",x"bf"),
   185 => (x"88",x"c1",x"48",x"87"),
   186 => (x"58",x"c9",x"ed",x"c2"),
   187 => (x"c1",x"87",x"ce",x"c0"),
   188 => (x"6a",x"4a",x"a5",x"d8"),
   189 => (x"87",x"c5",x"c0",x"02"),
   190 => (x"73",x"49",x"ff",x"4b"),
   191 => (x"48",x"a6",x"c4",x"0f"),
   192 => (x"49",x"74",x"78",x"c1"),
   193 => (x"c0",x"05",x"99",x"c4"),
   194 => (x"f2",x"c3",x"87",x"ce"),
   195 => (x"87",x"f5",x"e0",x"49"),
   196 => (x"99",x"c2",x"49",x"70"),
   197 => (x"87",x"ec",x"c0",x"02"),
   198 => (x"bf",x"c5",x"ed",x"c2"),
   199 => (x"b7",x"c7",x"48",x"7e"),
   200 => (x"cb",x"c0",x"03",x"a8"),
   201 => (x"c1",x"48",x"6e",x"87"),
   202 => (x"c9",x"ed",x"c2",x"80"),
   203 => (x"87",x"cf",x"c0",x"58"),
   204 => (x"7e",x"a5",x"d8",x"c1"),
   205 => (x"c0",x"02",x"bf",x"6e"),
   206 => (x"fe",x"4b",x"87",x"c5"),
   207 => (x"c4",x"0f",x"73",x"49"),
   208 => (x"78",x"c1",x"48",x"a6"),
   209 => (x"ff",x"49",x"fd",x"c3"),
   210 => (x"70",x"87",x"fa",x"df"),
   211 => (x"02",x"99",x"c2",x"49"),
   212 => (x"c2",x"87",x"e5",x"c0"),
   213 => (x"02",x"bf",x"c5",x"ed"),
   214 => (x"c2",x"87",x"c9",x"c0"),
   215 => (x"c0",x"48",x"c5",x"ed"),
   216 => (x"87",x"cf",x"c0",x"78"),
   217 => (x"7e",x"a5",x"d8",x"c1"),
   218 => (x"c0",x"02",x"bf",x"6e"),
   219 => (x"fd",x"4b",x"87",x"c5"),
   220 => (x"c4",x"0f",x"73",x"49"),
   221 => (x"78",x"c1",x"48",x"a6"),
   222 => (x"ff",x"49",x"fa",x"c3"),
   223 => (x"70",x"87",x"c6",x"df"),
   224 => (x"02",x"99",x"c2",x"49"),
   225 => (x"c2",x"87",x"e9",x"c0"),
   226 => (x"48",x"bf",x"c5",x"ed"),
   227 => (x"03",x"a8",x"b7",x"c7"),
   228 => (x"c2",x"87",x"c9",x"c0"),
   229 => (x"c7",x"48",x"c5",x"ed"),
   230 => (x"87",x"cf",x"c0",x"78"),
   231 => (x"7e",x"a5",x"d8",x"c1"),
   232 => (x"c0",x"02",x"bf",x"6e"),
   233 => (x"fc",x"4b",x"87",x"c5"),
   234 => (x"c4",x"0f",x"73",x"49"),
   235 => (x"78",x"c1",x"48",x"a6"),
   236 => (x"ed",x"c2",x"4b",x"c0"),
   237 => (x"50",x"c0",x"48",x"c0"),
   238 => (x"c4",x"49",x"ee",x"cb"),
   239 => (x"a6",x"cc",x"87",x"e5"),
   240 => (x"c0",x"ed",x"c2",x"58"),
   241 => (x"c1",x"05",x"bf",x"97"),
   242 => (x"49",x"74",x"87",x"de"),
   243 => (x"05",x"99",x"f0",x"c3"),
   244 => (x"c1",x"87",x"cd",x"c0"),
   245 => (x"dd",x"ff",x"49",x"da"),
   246 => (x"98",x"70",x"87",x"eb"),
   247 => (x"87",x"c8",x"c1",x"02"),
   248 => (x"bf",x"e8",x"4b",x"c1"),
   249 => (x"ff",x"c3",x"49",x"4c"),
   250 => (x"2c",x"b7",x"c8",x"99"),
   251 => (x"d3",x"c2",x"b4",x"71"),
   252 => (x"ff",x"49",x"bf",x"db"),
   253 => (x"c8",x"87",x"cb",x"d9"),
   254 => (x"f2",x"c3",x"49",x"66"),
   255 => (x"02",x"98",x"70",x"87"),
   256 => (x"c2",x"87",x"c6",x"c0"),
   257 => (x"c1",x"48",x"c0",x"ed"),
   258 => (x"c0",x"ed",x"c2",x"50"),
   259 => (x"c0",x"05",x"bf",x"97"),
   260 => (x"49",x"74",x"87",x"d6"),
   261 => (x"05",x"99",x"f0",x"c3"),
   262 => (x"c1",x"87",x"c5",x"ff"),
   263 => (x"dc",x"ff",x"49",x"da"),
   264 => (x"98",x"70",x"87",x"e3"),
   265 => (x"87",x"f8",x"fe",x"05"),
   266 => (x"c0",x"02",x"9b",x"73"),
   267 => (x"a6",x"c8",x"87",x"dc"),
   268 => (x"c5",x"ed",x"c2",x"48"),
   269 => (x"66",x"c8",x"78",x"bf"),
   270 => (x"75",x"91",x"cb",x"49"),
   271 => (x"bf",x"6e",x"7e",x"a1"),
   272 => (x"87",x"c6",x"c0",x"02"),
   273 => (x"49",x"66",x"c8",x"4b"),
   274 => (x"66",x"c4",x"0f",x"73"),
   275 => (x"87",x"c8",x"c0",x"02"),
   276 => (x"bf",x"c5",x"ed",x"c2"),
   277 => (x"87",x"e4",x"f1",x"49"),
   278 => (x"bf",x"df",x"d3",x"c2"),
   279 => (x"87",x"dd",x"c0",x"02"),
   280 => (x"87",x"cb",x"c2",x"49"),
   281 => (x"c0",x"02",x"98",x"70"),
   282 => (x"ed",x"c2",x"87",x"d3"),
   283 => (x"f1",x"49",x"bf",x"c5"),
   284 => (x"49",x"c0",x"87",x"ca"),
   285 => (x"c2",x"87",x"ea",x"f2"),
   286 => (x"c0",x"48",x"df",x"d3"),
   287 => (x"f2",x"8e",x"f4",x"78"),
   288 => (x"5e",x"0e",x"87",x"c4"),
   289 => (x"0e",x"5d",x"5c",x"5b"),
   290 => (x"c2",x"4c",x"71",x"1e"),
   291 => (x"49",x"bf",x"c1",x"ed"),
   292 => (x"4d",x"a1",x"cd",x"c1"),
   293 => (x"69",x"81",x"d1",x"c1"),
   294 => (x"02",x"9c",x"74",x"7e"),
   295 => (x"a5",x"c4",x"87",x"cf"),
   296 => (x"c2",x"7b",x"74",x"4b"),
   297 => (x"49",x"bf",x"c1",x"ed"),
   298 => (x"6e",x"87",x"e3",x"f1"),
   299 => (x"05",x"9c",x"74",x"7b"),
   300 => (x"4b",x"c0",x"87",x"c4"),
   301 => (x"4b",x"c1",x"87",x"c2"),
   302 => (x"e4",x"f1",x"49",x"73"),
   303 => (x"02",x"66",x"d4",x"87"),
   304 => (x"de",x"49",x"87",x"c7"),
   305 => (x"c2",x"4a",x"70",x"87"),
   306 => (x"c2",x"4a",x"c0",x"87"),
   307 => (x"26",x"5a",x"e3",x"d3"),
   308 => (x"00",x"87",x"f3",x"f0"),
   309 => (x"00",x"00",x"00",x"00"),
   310 => (x"00",x"00",x"00",x"00"),
   311 => (x"00",x"00",x"00",x"00"),
   312 => (x"1e",x"00",x"00",x"00"),
   313 => (x"c8",x"ff",x"4a",x"71"),
   314 => (x"a1",x"72",x"49",x"bf"),
   315 => (x"1e",x"4f",x"26",x"48"),
   316 => (x"89",x"bf",x"c8",x"ff"),
   317 => (x"c0",x"c0",x"c0",x"fe"),
   318 => (x"01",x"a9",x"c0",x"c0"),
   319 => (x"4a",x"c0",x"87",x"c4"),
   320 => (x"4a",x"c1",x"87",x"c2"),
   321 => (x"4f",x"26",x"48",x"72"),
   322 => (x"5c",x"5b",x"5e",x"0e"),
   323 => (x"4b",x"71",x"0e",x"5d"),
   324 => (x"d0",x"4c",x"d4",x"ff"),
   325 => (x"78",x"c0",x"48",x"66"),
   326 => (x"da",x"ff",x"49",x"d6"),
   327 => (x"ff",x"c3",x"87",x"df"),
   328 => (x"c3",x"49",x"6c",x"7c"),
   329 => (x"4d",x"71",x"99",x"ff"),
   330 => (x"99",x"f0",x"c3",x"49"),
   331 => (x"05",x"a9",x"e0",x"c1"),
   332 => (x"ff",x"c3",x"87",x"cb"),
   333 => (x"c3",x"48",x"6c",x"7c"),
   334 => (x"08",x"66",x"d0",x"98"),
   335 => (x"7c",x"ff",x"c3",x"78"),
   336 => (x"c8",x"49",x"4a",x"6c"),
   337 => (x"7c",x"ff",x"c3",x"31"),
   338 => (x"b2",x"71",x"4a",x"6c"),
   339 => (x"31",x"c8",x"49",x"72"),
   340 => (x"6c",x"7c",x"ff",x"c3"),
   341 => (x"72",x"b2",x"71",x"4a"),
   342 => (x"c3",x"31",x"c8",x"49"),
   343 => (x"4a",x"6c",x"7c",x"ff"),
   344 => (x"d0",x"ff",x"b2",x"71"),
   345 => (x"78",x"e0",x"c0",x"48"),
   346 => (x"c2",x"02",x"9b",x"73"),
   347 => (x"75",x"7b",x"72",x"87"),
   348 => (x"26",x"4d",x"26",x"48"),
   349 => (x"26",x"4b",x"26",x"4c"),
   350 => (x"4f",x"26",x"1e",x"4f"),
   351 => (x"5c",x"5b",x"5e",x"0e"),
   352 => (x"76",x"86",x"f8",x"0e"),
   353 => (x"49",x"a6",x"c8",x"1e"),
   354 => (x"c4",x"87",x"fd",x"fd"),
   355 => (x"6e",x"4b",x"70",x"86"),
   356 => (x"01",x"a8",x"c0",x"48"),
   357 => (x"73",x"87",x"f0",x"c2"),
   358 => (x"9a",x"f0",x"c3",x"4a"),
   359 => (x"02",x"aa",x"d0",x"c1"),
   360 => (x"e0",x"c1",x"87",x"c7"),
   361 => (x"de",x"c2",x"05",x"aa"),
   362 => (x"c8",x"49",x"73",x"87"),
   363 => (x"87",x"c3",x"02",x"99"),
   364 => (x"73",x"87",x"c6",x"ff"),
   365 => (x"c2",x"9c",x"c3",x"4c"),
   366 => (x"c2",x"c1",x"05",x"ac"),
   367 => (x"49",x"66",x"c4",x"87"),
   368 => (x"1e",x"71",x"31",x"c9"),
   369 => (x"d4",x"4a",x"66",x"c4"),
   370 => (x"c9",x"ed",x"c2",x"92"),
   371 => (x"fe",x"81",x"72",x"49"),
   372 => (x"d8",x"87",x"f4",x"cf"),
   373 => (x"e4",x"d7",x"ff",x"49"),
   374 => (x"1e",x"c0",x"c8",x"87"),
   375 => (x"49",x"f2",x"db",x"c2"),
   376 => (x"87",x"fa",x"eb",x"fd"),
   377 => (x"c0",x"48",x"d0",x"ff"),
   378 => (x"db",x"c2",x"78",x"e0"),
   379 => (x"66",x"cc",x"1e",x"f2"),
   380 => (x"c2",x"92",x"d4",x"4a"),
   381 => (x"72",x"49",x"c9",x"ed"),
   382 => (x"fc",x"cd",x"fe",x"81"),
   383 => (x"c1",x"86",x"cc",x"87"),
   384 => (x"c2",x"c1",x"05",x"ac"),
   385 => (x"49",x"66",x"c4",x"87"),
   386 => (x"1e",x"71",x"31",x"c9"),
   387 => (x"d4",x"4a",x"66",x"c4"),
   388 => (x"c9",x"ed",x"c2",x"92"),
   389 => (x"fe",x"81",x"72",x"49"),
   390 => (x"c2",x"87",x"ec",x"ce"),
   391 => (x"c8",x"1e",x"f2",x"db"),
   392 => (x"92",x"d4",x"4a",x"66"),
   393 => (x"49",x"c9",x"ed",x"c2"),
   394 => (x"cb",x"fe",x"81",x"72"),
   395 => (x"49",x"d7",x"87",x"fd"),
   396 => (x"87",x"c9",x"d6",x"ff"),
   397 => (x"c2",x"1e",x"c0",x"c8"),
   398 => (x"fd",x"49",x"f2",x"db"),
   399 => (x"cc",x"87",x"f8",x"e9"),
   400 => (x"48",x"d0",x"ff",x"86"),
   401 => (x"f8",x"78",x"e0",x"c0"),
   402 => (x"87",x"e7",x"fc",x"8e"),
   403 => (x"5c",x"5b",x"5e",x"0e"),
   404 => (x"4a",x"71",x"0e",x"5d"),
   405 => (x"d0",x"4c",x"d4",x"ff"),
   406 => (x"b7",x"c3",x"4d",x"66"),
   407 => (x"87",x"c5",x"06",x"ad"),
   408 => (x"e1",x"c1",x"48",x"c0"),
   409 => (x"75",x"1e",x"72",x"87"),
   410 => (x"c2",x"93",x"d4",x"4b"),
   411 => (x"73",x"83",x"c9",x"ed"),
   412 => (x"c4",x"c6",x"fe",x"49"),
   413 => (x"6b",x"83",x"c8",x"87"),
   414 => (x"48",x"d0",x"ff",x"4b"),
   415 => (x"dd",x"78",x"e1",x"c8"),
   416 => (x"c3",x"48",x"73",x"7c"),
   417 => (x"7c",x"70",x"98",x"ff"),
   418 => (x"b7",x"c8",x"49",x"73"),
   419 => (x"c3",x"48",x"71",x"29"),
   420 => (x"7c",x"70",x"98",x"ff"),
   421 => (x"b7",x"d0",x"49",x"73"),
   422 => (x"c3",x"48",x"71",x"29"),
   423 => (x"7c",x"70",x"98",x"ff"),
   424 => (x"b7",x"d8",x"48",x"73"),
   425 => (x"c0",x"7c",x"70",x"28"),
   426 => (x"7c",x"7c",x"7c",x"7c"),
   427 => (x"7c",x"7c",x"7c",x"7c"),
   428 => (x"7c",x"7c",x"7c",x"7c"),
   429 => (x"c0",x"48",x"d0",x"ff"),
   430 => (x"1e",x"75",x"78",x"e0"),
   431 => (x"d4",x"ff",x"49",x"dc"),
   432 => (x"86",x"c8",x"87",x"e0"),
   433 => (x"e8",x"fa",x"48",x"73"),
   434 => (x"e8",x"fa",x"48",x"87"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

